* BEGIN ANSOFT HEADER
* node 1    DC+:D1K
* node 2    DC+:D2K
* node 3    DC+:D3K
* node 4    DC+:D4K
* node 5    DC-:DC-GS-short-b
* node 6    DC-:Q1BW
* node 7    DC-:Q1S
* node 8    DC-:Q2BW
* node 9    DC-:Q2S
* node 10   DC-:Q3BW
* node 11   DC-:Q3S
* node 12   DC-:Q4BW
* node 13   DC-:Q4S
* node 14   DC-:RS1b
* node 15   DC-:RS2b
* node 16   DC-:RS3b
* node 17   DC-:RS4b
* node 18   G1:Q1G
* node 19   G2:Q2G
* node 20   G3:Q3G
* node 21   G4:Q4G
* node 22   GG:RG1a
* node 23   GG:RG2a
* node 24   GG:RG3a
* node 25   GG:RG4a
* node 26   GS:DC-GS-short-a
* node 27   GS:RS1a
* node 28   GS:RS2a
* node 29   GS:RS3a
* node 30   GS:RS4a
* node 31   OUT:D1A
* node 32   OUT:D2A
* node 33   OUT:D3A
* node 34   OUT:D4A
* node 35   OUT:Q1D
* node 36   OUT:Q2D
* node 37   OUT:Q3D
* node 38   OUT:Q4D
* node 39   DC+:DC+terminal
* node 40   DC-:DC-terminal
* node 41   G1:RG1b
* node 42   G2:RG2b
* node 43   G3:RG3b
* node 44   G4:RG4b
* node 45   GG:G-terminal
* node 46   GS:S-terminal
* node 47   OUT:OUT-terminal
*  Project: Quadraat
*   Design: Q3DDesign1
*   Format: Ansys Nexxim
*   Topckt: Quadraat
*  Creator: Ansys Electronics Desktop 2022.1.0
*     Date: Fri Nov 18 10:37:14 2022
* END ANSOFT HEADER

.subckt Quadraat 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24
+ 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42 43 44 45 46 47
X1 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29
+ 30 31 32 33 34 35 36 37 38 39 39 39 39 40 40 40 40 40 40 40 40 40 40 40 40 40
+ 41 42 43 44 45 45 45 45 46 46 46 46 46 47 47 47 47 47 47 47 47 Quadraat_series

.subckt Quadraat_series 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22
+ 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42 43 44 45 46 47 48
+ 49 50 51 52 53 54 55 56 57 58 59 60 61 62 63 64 65 66 67 68 69 70 71 72 73 74
+ 75 76
V1 1 77 dc 0.0
V2 2 78 dc 0.0
V3 3 79 dc 0.0
V4 4 80 dc 0.0
V5 5 81 dc 0.0
V6 6 82 dc 0.0
V7 7 83 dc 0.0
V8 8 84 dc 0.0
V9 9 85 dc 0.0
V10 10 86 dc 0.0
V11 11 87 dc 0.0
V12 12 88 dc 0.0
V13 13 89 dc 0.0
V14 14 90 dc 0.0
V15 15 91 dc 0.0
V16 16 92 dc 0.0
V17 17 93 dc 0.0
V18 18 94 dc 0.0
V19 19 95 dc 0.0
V20 20 96 dc 0.0
V21 21 97 dc 0.0
V22 22 98 dc 0.0
V23 23 99 dc 0.0
V24 24 100 dc 0.0
V25 25 101 dc 0.0
V26 26 102 dc 0.0
V27 27 103 dc 0.0
V28 28 104 dc 0.0
V29 29 105 dc 0.0
V30 30 106 dc 0.0
V31 31 107 dc 0.0
V32 32 108 dc 0.0
V33 33 109 dc 0.0
V34 34 110 dc 0.0
V35 35 111 dc 0.0
V36 36 112 dc 0.0
V37 37 113 dc 0.0
V38 38 114 dc 0.0
R1 77 115 0.00101526580168
R2 78 116 0.00096894723124
R3 79 117 0.000923668356411
R4 80 118 0.000878053277473
R5 81 119 0.000900223586849
R6 82 120 0.000984291031383
R7 83 121 0.00262485569584
R8 84 122 0.00106983569313
R9 85 123 0.00271365819285
R10 86 124 0.00115311636051
R11 87 125 0.00279287283507
R12 88 126 0.00123800637645
R13 89 127 0.00288202449098
R14 90 128 0.00659941879782
R15 91 129 0.00668981503575
R16 92 130 0.00678076942227
R17 93 131 0.00685916426004
R18 94 132 0.00365468664321
R19 95 133 0.00365086260863
R20 96 134 0.00366949603563
R21 97 135 0.00365804213476
R22 98 136 0.00540231001262
R23 99 137 0.00500049155772
R24 100 138 0.00459671364279
R25 101 139 0.00419503426918
R26 102 140 0.00466243404098
R27 103 141 0.00463192129081
R28 104 142 0.00423263467888
R29 105 143 0.00383687377396
R30 106 144 0.00344111216291
R31 107 145 0.00181620034651
R32 108 146 0.00194313930967
R33 109 147 0.00205958004544
R34 110 148 0.00218704021588
R35 111 149 0.000494520671913
R36 112 150 0.000449759089926
R37 113 151 0.000405068333812
R38 114 152 0.000361298438952
F1_2 115 77 V2 0.954109
F1_3 115 77 V3 0.909521
F1_4 115 77 V4 0.864677
F2_1 116 78 V1 0.999718
F2_3 116 78 V3 0.952999
F2_4 116 78 V4 0.906011
F3_1 117 79 V1 0.999715
F3_2 117 79 V2 0.999716
F3_4 117 79 V4 0.950425
F4_1 118 80 V1 0.999799
F4_2 118 80 V2 0.999799
F4_3 118 80 V3 0.9998
F5_6 119 81 V6 0.910453
F5_7 119 81 V7 0.910453
F5_8 119 81 V8 0.910447
F5_9 119 81 V9 0.910447
F5_10 119 81 V10 0.910447
F5_11 119 81 V11 0.910447
F5_12 119 81 V12 0.910447
F5_13 119 81 V13 0.910447
F5_14 119 81 V14 0.910453
F5_15 119 81 V15 0.910447
F5_16 119 81 V16 0.910447
F5_17 119 81 V17 0.910447
F6_5 120 82 V5 0.832692
F6_7 120 82 V7 0.997817
F6_8 120 82 V8 0.985357
F6_9 120 82 V9 0.985361
F6_10 120 82 V10 0.985214
F6_11 120 82 V11 0.985214
F6_12 120 82 V12 0.985212
F6_13 120 82 V13 0.985212
F6_14 120 82 V14 0.997817
F6_15 120 82 V15 0.985361
F6_16 120 82 V16 0.985214
F6_17 120 82 V17 0.985212
F7_5 121 83 V5 0.31225
F7_6 121 83 V6 0.37417
F7_8 121 83 V8 0.369521
F7_9 121 83 V9 0.369523
F7_10 121 83 V10 0.369464
F7_11 121 83 V11 0.369464
F7_12 121 83 V12 0.369463
F7_13 121 83 V13 0.369463
F7_14 121 83 V14 0.999996
F7_15 121 83 V15 0.369523
F7_16 121 83 V16 0.369464
F7_17 121 83 V17 0.369463
F8_5 122 84 V5 0.766104
F8_6 122 84 V6 0.906567
F8_7 122 84 V7 0.906625
F8_9 122 84 V9 0.995712
F8_10 122 84 V10 0.982855
F8_11 122 84 V11 0.98286
F8_12 122 84 V12 0.982704
F8_13 122 84 V13 0.982704
F8_14 122 84 V14 0.906625
F8_15 122 84 V15 0.995712
F8_16 122 84 V16 0.98286
F8_17 122 84 V17 0.982704
F9_5 123 85 V5 0.30203
F9_6 123 85 V6 0.357408
F9_7 123 85 V7 0.357431
F9_8 123 85 V8 0.392551
F9_10 123 85 V10 0.387586
F9_11 123 85 V11 0.387588
F9_12 123 85 V12 0.387523
F9_13 123 85 V13 0.387523
F9_14 123 85 V14 0.357431
F9_15 123 85 V15 1
F9_16 123 85 V16 0.387588
F9_17 123 85 V17 0.387523
F10_5 124 86 V5 0.710774
F10_6 124 86 V6 0.840971
F10_7 124 86 V7 0.841016
F10_8 124 86 V8 0.911871
F10_9 124 86 V9 0.912116
F10_11 124 86 V11 0.994761
F10_12 124 86 V12 0.982243
F10_13 124 86 V13 0.98225
F10_14 124 86 V14 0.841016
F10_15 124 86 V15 0.912116
F10_16 124 86 V16 0.994761
F10_17 124 86 V17 0.98225
F11_5 125 87 V5 0.293463
F11_6 125 87 V6 0.347218
F11_7 125 87 V7 0.347237
F11_8 125 87 V8 0.376494
F11_9 125 87 V9 0.376595
F11_10 125 87 V10 0.410715
F11_12 125 87 V12 0.405623
F11_13 125 87 V13 0.405626
F11_14 125 87 V14 0.347237
F11_15 125 87 V15 0.376595
F11_16 125 87 V16 0.999996
F11_17 125 87 V17 0.405626
F12_5 126 88 V5 0.662037
F12_6 126 88 V6 0.783304
F12_7 126 88 V7 0.783346
F12_8 126 88 V8 0.849214
F12_9 126 88 V9 0.849435
F12_10 126 88 V10 0.914891
F12_11 126 88 V11 0.915062
F12_13 126 88 V13 0.996014
F12_14 126 88 V14 0.783346
F12_15 126 88 V15 0.849435
F12_16 126 88 V16 0.915062
F12_17 126 88 V17 0.996014
F13_5 127 89 V5 0.284385
F13_6 127 89 V6 0.336477
F13_7 127 89 V7 0.336495
F13_8 127 89 V8 0.364789
F13_9 127 89 V9 0.364884
F13_10 127 89 V10 0.393005
F13_11 127 89 V11 0.393078
F13_12 127 89 V12 0.427849
F13_14 127 89 V14 0.336495
F13_15 127 89 V15 0.364884
F13_16 127 89 V16 0.393078
F13_17 127 89 V17 1
F14_5 128 90 V5 0.124194
F14_6 128 90 V6 0.148823
F14_7 128 90 V7 0.397739
F14_8 128 90 V8 0.146974
F14_9 128 90 V9 0.146974
F14_10 128 90 V10 0.146951
F14_11 128 90 V11 0.146951
F14_12 128 90 V12 0.14695
F14_13 128 90 V13 0.14695
F14_15 128 90 V15 0.146974
F14_16 128 90 V16 0.146951
F14_17 128 90 V17 0.14695
F15_5 129 91 V5 0.122515
F15_6 129 91 V6 0.144979
F15_7 129 91 V7 0.144988
F15_8 129 91 V8 0.159234
F15_9 129 91 V9 0.40564
F15_10 129 91 V10 0.157221
F15_11 129 91 V11 0.157221
F15_12 129 91 V12 0.157195
F15_13 129 91 V13 0.157195
F15_14 129 91 V14 0.144988
F15_16 129 91 V16 0.157221
F15_17 129 91 V17 0.157195
F16_5 130 92 V5 0.120872
F16_6 130 92 V6 0.143013
F16_7 130 92 V7 0.143021
F16_8 130 92 V8 0.155071
F16_9 130 92 V9 0.155113
F16_10 130 92 V10 0.169166
F16_11 130 92 V11 0.41188
F16_12 130 92 V12 0.167068
F16_13 130 92 V13 0.16707
F16_14 130 92 V14 0.143021
F16_15 130 92 V15 0.155113
F16_17 130 92 V17 0.16707
F17_5 131 93 V5 0.119491
F17_6 131 93 V6 0.141378
F17_7 131 93 V7 0.141386
F17_8 131 93 V8 0.153274
F17_9 131 93 V9 0.153314
F17_10 131 93 V10 0.165129
F17_11 131 93 V11 0.16516
F17_12 131 93 V12 0.17977
F17_13 131 93 V13 0.420171
F17_14 131 93 V14 0.141386
F17_15 131 93 V15 0.153314
F17_16 131 93 V16 0.16516
F22_23 136 98 V23 0.925604
F22_24 136 98 V24 0.850861
F22_25 136 98 V25 0.776505
F23_22 137 99 V22 0.999982
F23_24 137 99 V24 0.919233
F23_25 137 99 V25 0.838902
F24_22 138 100 V22 0.999979
F24_23 138 100 V23 0.999979
F24_25 138 100 V25 0.912591
F25_22 139 101 V22 0.999973
F25_23 139 101 V23 0.999973
F25_24 139 101 V24 0.999973
F26_27 140 102 V27 0.993431
F26_28 140 102 V28 0.907795
F26_29 140 102 V29 0.822922
F26_30 140 102 V30 0.738015
F27_26 141 103 V26 0.999976
F27_28 141 103 V28 0.913775
F27_29 141 103 V29 0.828343
F27_30 141 103 V30 0.742877
F28_26 142 104 V26 0.999977
F28_27 142 104 V27 0.999977
F28_29 142 104 V29 0.906485
F28_30 142 104 V30 0.812956
F29_26 143 105 V26 0.999986
F29_27 143 105 V27 0.999986
F29_28 143 105 V28 0.999986
F29_30 143 105 V30 0.89681
F30_26 144 106 V26 0.999952
F30_27 144 106 V27 0.999952
F30_28 144 106 V28 0.999952
F30_29 144 106 V29 0.999952
F31_32 145 107 V32 0.105261
F31_33 145 107 V33 0.105197
F31_34 145 107 V34 0.105207
F31_35 145 107 V35 0.0551517
F31_36 145 107 V36 0.0551517
F31_37 145 107 V37 0.0551517
F31_38 145 107 V38 0.0551517
F32_31 146 108 V31 0.0983851
F32_33 146 108 V33 0.161642
F32_34 146 108 V34 0.161575
F32_35 146 108 V35 0.0515158
F32_36 146 108 V36 0.0515158
F32_37 146 108 V37 0.0515158
F32_38 146 108 V38 0.0515158
F33_31 147 109 V31 0.092766
F33_32 147 109 V32 0.152504
F33_34 147 109 V34 0.211903
F33_35 147 109 V35 0.048604
F33_36 147 109 V36 0.048604
F33_37 147 109 V37 0.048604
F33_38 147 109 V38 0.048604
F34_31 148 110 V31 0.0873675
F34_32 148 110 V32 0.143556
F34_33 148 110 V33 0.199553
F34_35 148 110 V35 0.0457712
F34_36 148 110 V36 0.0457712
F34_37 148 110 V37 0.0457712
F34_38 148 110 V38 0.0457712
F35_31 149 111 V31 0.202553
F35_32 149 111 V32 0.202423
F35_33 149 111 V33 0.202426
F35_34 149 111 V34 0.202425
F35_36 149 111 V36 0.906734
F35_37 149 111 V37 0.816251
F35_38 149 111 V38 0.727012
F36_31 150 112 V31 0.222711
F36_32 150 112 V32 0.222569
F36_33 150 112 V33 0.222572
F36_34 150 112 V34 0.222571
F36_35 150 112 V35 0.996975
F36_37 150 112 V37 0.897498
F36_38 150 112 V38 0.799367
F37_31 151 113 V31 0.247283
F37_32 151 113 V32 0.247125
F37_33 151 113 V33 0.247128
F37_34 151 113 V34 0.247128
F37_35 151 113 V35 0.996506
F37_36 151 113 V36 0.996518
F37_38 151 113 V38 0.887573
F38_31 152 114 V31 0.27724
F38_32 152 114 V32 0.277063
F38_33 152 114 V33 0.277067
F38_34 152 114 V34 0.277066
F38_35 152 114 V35 0.995084
F38_36 152 114 V36 0.995084
F38_37 152 114 V37 0.9951
L1 115 39 9.87367044122e-09
L2 116 40 9.19764894195e-09
L3 117 41 8.47567530558e-09
L4 118 42 7.6793692027e-09
L5 119 43 7.25832700673e-09
L6 120 44 8.82690206486e-09
L7 121 45 1.08383687852e-08
L8 122 46 1.01626865639e-08
L9 123 47 1.23037878625e-08
L10 124 48 1.14238192044e-08
L11 125 49 1.36185759059e-08
L12 126 50 1.27138850898e-08
L13 127 51 1.49353915992e-08
L14 128 52 1.46478208018e-08
L15 129 53 1.62681093797e-08
L16 130 54 1.76170625661e-08
L17 131 55 1.89567082538e-08
L18 132 56 3.64633389566e-09
L19 133 57 3.64639708022e-09
L20 134 58 3.64845333175e-09
L21 135 59 3.66795804795e-09
L22 136 60 1.77593168857e-08
L23 137 61 1.60630849818e-08
L24 138 62 1.43086712787e-08
L25 139 63 1.24681750846e-08
L26 140 64 1.73032098316e-08
L27 141 65 1.70600690675e-08
L28 142 66 1.52336477298e-08
L29 143 67 1.33971096208e-08
L30 144 68 1.15006159027e-08
L31 145 69 4.33215568887e-09
L32 146 70 5.85684164769e-09
L33 147 71 7.40679037617e-09
L34 148 72 9.00157175731e-09
L35 149 73 6.74819853873e-09
L36 150 74 6.16048290132e-09
L37 151 75 5.70820968729e-09
L38 152 76 5.4437915387e-09
K1_2 L1 L2 0.970265
K1_3 L1 L3 0.936903
K1_4 L1 L4 0.901667
K1_5 L1 L5 0.14395
K1_6 L1 L6 0.133787
K1_7 L1 L7 0.126822
K1_8 L1 L8 0.158461
K1_9 L1 L9 0.143597
K1_10 L1 L10 0.174303
K1_11 L1 L11 0.155077
K1_12 L1 L12 0.18062
K1_13 L1 L13 0.160439
K1_14 L1 L14 0.109417
K1_15 L1 L15 0.124032
K1_16 L1 L16 0.13441
K1_17 L1 L17 0.139895
K1_18 L1 L18 -0.00735334
K1_19 L1 L19 -0.00370259
K1_20 L1 L20 -0.000660246
K1_21 L1 L21 0.00139338
K1_22 L1 L22 -0.00905795
K1_23 L1 L23 0.0003557
K1_24 L1 L24 0.00927632
K1_25 L1 L25 0.0166995
K1_26 L1 L26 -0.0107955
K1_27 L1 L27 -0.00764916
K1_28 L1 L28 0.00202833
K1_29 L1 L29 0.0116461
K1_30 L1 L30 0.0203891
K1_31 L1 L31 -0.0225915
K1_32 L1 L32 -0.0716663
K1_33 L1 L33 -0.120122
K1_34 L1 L34 -0.168178
K1_35 L1 L35 -0.107624
K1_36 L1 L36 -0.0887928
K1_37 L1 L37 -0.071848
K1_38 L1 L38 -0.058632
K2_3 L2 L3 0.967193
K2_4 L2 L4 0.93116
K2_5 L2 L5 0.14505
K2_6 L2 L6 0.137296
K2_7 L2 L7 0.128482
K2_8 L2 L8 0.159709
K2_9 L2 L9 0.143281
K2_10 L2 L10 0.169345
K2_11 L2 L11 0.150789
K2_12 L2 L12 0.169548
K2_13 L2 L13 0.152268
K2_14 L2 L14 0.110395
K2_15 L2 L15 0.123474
K2_16 L2 L16 0.130822
K2_17 L2 L17 0.133329
K2_18 L2 L18 -0.006207
K2_19 L2 L19 -0.00251799
K2_20 L2 L20 -0.000156415
K2_21 L2 L21 0.000842066
K2_22 L2 L22 -0.00394832
K2_23 L2 L23 0.00463581
K2_24 L2 L24 0.0121302
K2_25 L2 L25 0.0181327
K2_26 L2 L26 -0.00591018
K2_27 L2 L27 -0.0029084
K2_28 L2 L28 0.00610672
K2_29 L2 L29 0.014484
K2_30 L2 L30 0.0217939
K2_31 L2 L31 -0.0107795
K2_32 L2 L32 -0.0241766
K2_33 L2 L33 -0.0728395
K2_34 L2 L34 -0.126254
K2_35 L2 L35 -0.0776954
K2_36 L2 L36 -0.0595913
K2_37 L2 L37 -0.0456458
K2_38 L2 L38 -0.0362002
K3_4 L3 L4 0.96443
K3_5 L3 L5 0.144636
K3_6 L3 L6 0.140378
K3_7 L3 L7 0.128949
K3_8 L3 L8 0.156405
K3_9 L3 L9 0.139604
K3_10 L3 L10 0.158671
K3_11 L3 L11 0.142494
K3_12 L3 L12 0.156125
K3_13 L3 L13 0.141675
K3_14 L3 L14 0.110167
K3_15 L3 L15 0.12016
K3_16 L3 L16 0.12396
K3_17 L3 L17 0.124575
K3_18 L3 L18 -0.00449987
K3_19 L3 L19 -0.00142025
K3_20 L3 L20 -9.13689e-05
K3_21 L3 L21 0.000249282
K3_22 L3 L22 0.00171853
K3_23 L3 L23 0.00893526
K3_24 L3 L24 0.0147912
K3_25 L3 L25 0.0195932
K3_26 L3 L26 -0.000139949
K3_27 L3 L27 0.00258043
K3_28 L3 L28 0.0104642
K3_29 L3 L29 0.0173066
K3_30 L3 L30 0.0232795
K3_31 L3 L31 -0.00650316
K3_32 L3 L32 -0.0126487
K3_33 L3 L33 -0.0278154
K3_34 L3 L34 -0.0807978
K3_35 L3 L35 -0.0514326
K3_36 L3 L36 -0.0361212
K3_37 L3 L37 -0.0261546
K3_38 L3 L38 -0.0195083
K4_5 L4 L5 0.142137
K4_6 L4 L6 0.139897
K4_7 L4 L7 0.126648
K4_8 L4 L8 0.147258
K4_9 L4 L9 0.132114
K4_10 L4 L10 0.145918
K4_11 L4 L11 0.13222
K4_12 L4 L12 0.142512
K4_13 L4 L13 0.13031
K4_14 L4 L14 0.107629
K4_15 L4 L15 0.11381
K4_16 L4 L16 0.115371
K4_17 L4 L17 0.114951
K4_18 L4 L18 -0.00272156
K4_19 L4 L19 -0.000802859
K4_20 L4 L20 -0.000192835
K4_21 L4 L21 -0.00014011
K4_22 L4 L22 0.00710152
K4_23 L4 L23 0.0127849
K4_24 L4 L24 0.0173345
K4_25 L4 L25 0.0213244
K4_26 L4 L26 0.00574667
K4_27 L4 L27 0.00802923
K4_28 L4 L28 0.0145407
K4_29 L4 L29 0.0200233
K4_30 L4 L30 0.0250151
K4_31 L4 L31 -0.00392942
K4_32 L4 L32 -0.00923552
K4_33 L4 L33 -0.0174833
K4_34 L4 L34 -0.0387776
K4_35 L4 L35 -0.0319077
K4_36 L4 L36 -0.0205692
K4_37 L4 L37 -0.013603
K4_38 L4 L38 -0.00870115
K5_6 L5 L6 0.82731
K5_7 L5 L7 0.755272
K5_8 L5 L8 0.788333
K5_9 L5 L9 0.721269
K5_10 L5 L10 0.749934
K5_11 L5 L11 0.68998
K5_12 L5 L12 0.71438
K5_13 L5 L13 0.66128
K5_14 L5 L14 0.654407
K5_15 L5 L15 0.629948
K5_16 L5 L16 0.608114
K5_17 L5 L17 0.587885
K5_18 L5 L18 -0.0135829
K5_19 L5 L19 -0.0054443
K5_20 L5 L20 -0.00314797
K5_21 L5 L21 -0.00268855
K5_22 L5 L22 0.016001
K5_23 L5 L23 0.0190197
K5_24 L5 L24 0.0214656
K5_25 L5 L25 0.0243999
K5_26 L5 L26 0.00938397
K5_27 L5 L27 0.0172656
K5_28 L5 L28 0.0225827
K5_29 L5 L29 0.025946
K5_30 L5 L30 0.0298261
K5_31 L5 L31 -0.00145199
K5_32 L5 L32 -0.00935557
K5_33 L5 L33 -0.0193154
K5_34 L5 L34 -0.0334975
K5_35 L5 L35 -0.00388633
K5_36 L5 L36 0.00923555
K5_37 L5 L37 0.0143967
K5_38 L5 L38 0.0178628
K6_7 L6 L7 0.886092
K6_8 L6 L8 0.931752
K6_9 L6 L9 0.839341
K6_10 L6 L10 0.881283
K6_11 L6 L11 0.803127
K6_12 L6 L12 0.838377
K6_13 L6 L13 0.770688
K6_14 L6 L14 0.746076
K6_15 L6 L15 0.723956
K6_16 L6 L16 0.703226
K6_17 L6 L17 0.682134
K6_18 L6 L18 0.00829287
K6_19 L6 L19 0.00435395
K6_20 L6 L20 0.00248266
K6_21 L6 L21 0.00174303
K6_22 L6 L22 -0.00112953
K6_23 L6 L23 0.0128886
K6_24 L6 L24 0.0202361
K6_25 L6 L25 0.0253773
K6_26 L6 L26 -0.017886
K6_27 L6 L27 -0.00693397
K6_28 L6 L28 0.0123378
K6_29 L6 L29 0.0226019
K6_30 L6 L30 0.0296326
K6_31 L6 L31 -0.00486769
K6_32 L6 L32 -0.00643474
K6_33 L6 L33 -0.00952872
K6_34 L6 L34 -0.0221113
K6_35 L6 L35 -0.0551571
K6_36 L6 L36 -0.0352652
K6_37 L6 L37 -0.0277414
K6_38 L6 L38 -0.0227776
K7_8 L7 L8 0.827109
K7_9 L7 L9 0.754694
K7_10 L7 L10 0.783036
K7_11 L7 L11 0.717596
K7_12 L7 L12 0.745027
K7_13 L7 L13 0.68744
K7_14 L7 L14 0.848115
K7_15 L7 L15 0.654941
K7_16 L7 L16 0.630374
K7_17 L7 L17 0.609817
K7_18 L7 L18 0.00463477
K7_19 L7 L19 -0.00084867
K7_20 L7 L20 -0.000598465
K7_21 L7 L21 -0.000711558
K7_22 L7 L22 0.00202129
K7_23 L7 L23 0.0123838
K7_24 L7 L24 0.0173168
K7_25 L7 L25 0.0210302
K7_26 L7 L26 -0.0128086
K7_27 L7 L27 -0.00299247
K7_28 L7 L28 0.012826
K7_29 L7 L29 0.0202427
K7_30 L7 L30 0.0254284
K7_31 L7 L31 -0.00316487
K7_32 L7 L32 -0.00851013
K7_33 L7 L33 -0.0160081
K7_34 L7 L34 -0.0300706
K7_35 L7 L35 -0.0209258
K7_36 L7 L36 -0.00796868
K7_37 L7 L37 -0.00294092
K7_38 L7 L38 0.000789515
K8_9 L8 L9 0.900752
K8_10 L8 L10 0.940065
K8_11 L8 L11 0.856743
K8_12 L8 L12 0.893063
K8_13 L8 L13 0.821434
K8_14 L8 L14 0.697801
K8_15 L8 L15 0.775933
K8_16 L8 L16 0.749363
K8_17 L8 L17 0.726935
K8_18 L8 L18 0.00108608
K8_19 L8 L19 0.00319461
K8_20 L8 L20 0.00258536
K8_21 L8 L21 0.00141514
K8_22 L8 L22 -0.0173696
K8_23 L8 L23 0.00459387
K8_24 L8 L24 0.01554
K8_25 L8 L25 0.0218034
K8_26 L8 L26 -0.0348619
K8_27 L8 L27 -0.0230364
K8_28 L8 L28 0.00229341
K8_29 L8 L29 0.0172446
K8_30 L8 L30 0.0261846
K8_31 L8 L31 -0.00563844
K8_32 L8 L32 -0.0127947
K8_33 L8 L33 -0.03088
K8_34 L8 L34 -0.0613806
K8_35 L8 L35 -0.0866068
K8_36 L8 L36 -0.0360457
K8_37 L8 L37 -0.0214046
K8_38 L8 L38 -0.0152308
K9_10 L9 L10 0.848116
K9_11 L9 L11 0.781323
K9_12 L9 L12 0.806436
K9_13 L9 L13 0.745304
K9_14 L9 L14 0.640028
K9_15 L9 L15 0.864394
K9_16 L9 L16 0.686812
K9_17 L9 L17 0.661466
K9_18 L9 L18 -0.00596438
K9_19 L9 L19 0.00101936
K9_20 L9 L20 -0.00204399
K9_21 L9 L21 -0.00174952
K9_22 L9 L22 -0.0156819
K9_23 L9 L23 0.00513014
K9_24 L9 L24 0.0134036
K9_25 L9 L25 0.0179413
K9_26 L9 L26 -0.0317973
K9_27 L9 L27 -0.0208242
K9_28 L9 L28 0.00307386
K9_29 L9 L29 0.0157945
K9_30 L9 L30 0.0226444
K9_31 L9 L31 -0.00437612
K9_32 L9 L32 -0.0150427
K9_33 L9 L33 -0.0324847
K9_34 L9 L34 -0.0574012
K9_35 L9 L35 -0.0534281
K9_36 L9 L36 -0.00127903
K9_37 L9 L37 0.00767316
K9_38 L9 L38 0.0120259
K10_11 L10 L11 0.910807
K10_12 L10 L12 0.945318
K10_13 L10 L13 0.869307
K10_14 L10 L14 0.661449
K10_15 L10 L15 0.731627
K10_16 L10 L16 0.795346
K10_17 L10 L17 0.768334
K10_18 L10 L18 -0.00213711
K10_19 L10 L19 -0.00278293
K10_20 L10 L20 0.00182741
K10_21 L10 L21 0.00173449
K10_22 L10 L22 -0.0359149
K10_23 L10 L23 -0.0108758
K10_24 L10 L24 0.00825866
K10_25 L10 L25 0.0182637
K10_26 L10 L26 -0.0515334
K10_27 L10 L27 -0.0398571
K10_28 L10 L28 -0.0127635
K10_29 L10 L29 0.00863681
K10_30 L10 L30 0.0224831
K10_31 L10 L31 -0.00799744
K10_32 L10 L32 -0.0333816
K10_33 L10 L33 -0.0677216
K10_34 L10 L34 -0.100073
K10_35 L10 L35 -0.113978
K10_36 L10 L36 -0.0606185
K10_37 L10 L37 -0.0150925
K10_38 L10 L38 -0.00145485
K11_12 L11 L12 0.862473
K11_13 L11 L13 0.801188
K11_14 L11 L14 0.607941
K11_15 L11 L15 0.676802
K11_16 L11 L16 0.875545
K11_17 L11 L17 0.711433
K11_18 L11 L18 -0.0054702
K11_19 L11 L19 -0.00907142
K11_20 L11 L20 -0.000154476
K11_21 L11 L21 -0.00343061
K11_22 L11 L22 -0.036475
K11_23 L11 L23 -0.0123519
K11_24 L11 L24 0.00641758
K11_25 L11 L25 0.014422
K11_26 L11 L26 -0.0505749
K11_27 L11 L27 -0.0397327
K11_28 L11 L28 -0.0140058
K11_29 L11 L29 0.00690215
K11_30 L11 L30 0.019233
K11_31 L11 L31 -0.00718839
K11_32 L11 L32 -0.0298975
K11_33 L11 L33 -0.0576984
K11_34 L11 L34 -0.0850395
K11_35 L11 L35 -0.0762434
K11_36 L11 L36 -0.0240492
K11_37 L11 L37 0.024465
K11_38 L11 L38 0.0330402
K12_13 L12 L13 0.91859
K12_14 L12 L14 0.629571
K12_15 L12 L15 0.696407
K12_16 L12 L16 0.753973
K12_17 L12 L17 0.810076
K12_18 L12 L18 -0.0031359
K12_19 L12 L19 -0.00561234
K12_20 L12 L20 -0.00364753
K12_21 L12 L21 0.00187572
K12_22 L12 L22 -0.0521028
K12_23 L12 L23 -0.0274641
K12_24 L12 L24 -0.0049946
K12_25 L12 L25 0.0132991
K12_26 L12 L26 -0.0645837
K12_27 L12 L27 -0.053333
K12_28 L12 L28 -0.0269137
K12_29 L12 L29 -0.00336745
K12_30 L12 L30 0.0171919
K12_31 L12 L31 -0.0225916
K12_32 L12 L32 -0.0638292
K12_33 L12 L33 -0.0988415
K12_34 L12 L34 -0.128485
K12_35 L12 L35 -0.126683
K12_36 L12 L36 -0.0757063
K12_37 L12 L37 -0.0259083
K12_38 L12 L38 0.0202511
K13_14 L13 L14 0.582105
K13_15 L13 L15 0.645203
K13_16 L13 L16 0.703126
K13_17 L13 L17 0.884632
K13_18 L13 L18 -0.00517237
K13_19 L13 L19 -0.00870134
K13_20 L13 L20 -0.0101884
K13_21 L13 L21 -0.00210931
K13_22 L13 L22 -0.0554974
K13_23 L13 L23 -0.032173
K13_24 L13 L24 -0.00998574
K13_25 L13 L25 0.00875778
K13_26 L13 L26 -0.0659098
K13_27 L13 L27 -0.0554577
K13_28 L13 L28 -0.0306376
K13_29 L13 L29 -0.00770233
K13_30 L13 L30 0.0131403
K13_31 L13 L31 -0.0163263
K13_32 L13 L32 -0.0495473
K13_33 L13 L33 -0.0793289
K13_34 L13 L34 -0.105841
K13_35 L13 L35 -0.075015
K13_36 L13 L36 -0.0247952
K13_37 L13 L37 0.0254043
K13_38 L13 L38 0.0752104
K14_15 L14 L15 0.561826
K14_16 L14 L16 0.535772
K14_17 L14 L17 0.517269
K14_18 L14 L18 -0.1177
K14_19 L14 L19 -0.00798041
K14_20 L14 L20 -0.00288754
K14_21 L14 L21 -0.00206654
K14_22 L14 L22 0.00451924
K14_23 L14 L23 0.0105951
K14_24 L14 L24 0.0136814
K14_25 L14 L25 0.0163259
K14_26 L14 L26 -0.00804399
K14_27 L14 L27 0.00113472
K14_28 L14 L28 0.0120252
K14_29 L14 L29 0.0166566
K14_30 L14 L30 0.020317
K14_31 L14 L31 -0.00202964
K14_32 L14 L32 -0.00773922
K14_33 L14 L33 -0.0152904
K14_34 L14 L34 -0.0280577
K14_35 L14 L35 -0.012227
K14_36 L14 L36 0.00157833
K14_37 L14 L37 0.00624103
K14_38 L14 L38 0.00936072
K15_16 L15 L16 0.600658
K15_17 L15 L17 0.574237
K15_18 L15 L18 -0.0216569
K15_19 L15 L19 -0.114714
K15_20 L15 L20 -0.00870064
K15_21 L15 L21 -0.00396907
K15_22 L15 L22 -0.0122236
K15_23 L15 L23 0.00614849
K15_24 L15 L24 0.0108449
K15_25 L15 L25 0.013858
K15_26 L15 L26 -0.0268659
K15_27 L15 L27 -0.0170162
K15_28 L15 L28 0.00517918
K15_29 L15 L29 0.0138992
K15_30 L15 L30 0.0183643
K15_31 L15 L31 -0.00320215
K15_32 L15 L32 -0.0131974
K15_33 L15 L33 -0.0285126
K15_34 L15 L34 -0.0497086
K15_35 L15 L35 -0.0357659
K15_36 L15 L36 0.00459761
K15_37 L15 L37 0.0154626
K15_38 L15 L38 0.0197781
K16_17 L16 L17 0.629859
K16_18 L16 L18 -0.00826989
K16_19 L16 L19 -0.0237401
K16_20 L16 L20 -0.1113
K16_21 L16 L21 -0.0102122
K16_22 L16 L22 -0.0336526
K16_23 L16 L23 -0.0113257
K16_24 L16 L24 0.00535224
K16_25 L16 L25 0.00994161
K16_26 L16 L26 -0.0464993
K16_27 L16 L27 -0.0368762
K16_28 L16 L28 -0.0134029
K16_29 L16 L29 0.00654374
K16_30 L16 L30 0.0151172
K16_31 L16 L31 -0.00548485
K16_32 L16 L32 -0.0250509
K16_33 L16 L33 -0.0486377
K16_34 L16 L34 -0.0720561
K16_35 L16 L35 -0.0549177
K16_36 L16 L36 -0.00925345
K16_37 L16 L37 0.0286894
K16_38 L16 L38 0.0394086
K17_18 L17 L18 -0.00623931
K17_19 L17 L19 -0.011247
K17_20 L17 L20 -0.0247241
K17_21 L17 L21 -0.110407
K17_22 L17 L22 -0.0569155
K17_23 L17 L23 -0.0360738
K17_24 L17 L24 -0.01537
K17_25 L17 L25 0.00137989
K17_26 L17 L26 -0.0656192
K17_27 L17 L27 -0.0563411
K17_28 L17 L28 -0.0342762
K17_29 L17 L29 -0.0131426
K17_30 L17 L30 0.00710133
K17_31 L17 L31 -0.0125081
K17_32 L17 L32 -0.0405942
K17_33 L17 L33 -0.0661198
K17_34 L17 L34 -0.0892538
K17_35 L17 L35 -0.0516945
K17_36 L17 L36 -0.00629667
K17_37 L17 L37 0.0382732
K17_38 L17 L38 0.0776629
K18_19 L18 L19 0.0192088
K18_20 L18 L20 0.0050378
K18_21 L18 L21 0.00295247
K18_22 L18 L22 0.00164007
K18_23 L18 L23 0.00085139
K18_24 L18 L24 0.0022421
K18_25 L18 L25 0.00284886
K18_26 L18 L26 0.004834
K18_27 L18 L27 0.00270496
K18_28 L18 L28 -0.000594673
K18_29 L18 L29 0.001118
K18_30 L18 L30 0.00199214
K18_31 L18 L31 -0.000414999
K18_32 L18 L32 0.002639
K18_33 L18 L33 0.0058515
K18_34 L18 L34 0.0084245
K18_35 L18 L35 0.0020719
K18_36 L18 L36 -0.0129061
K18_37 L18 L37 -0.0156949
K18_38 L18 L38 -0.0164188
K19_20 L19 L20 0.019316
K19_21 L19 L21 0.00574582
K19_22 L19 L22 0.0114115
K19_23 L19 L23 0.00362122
K19_24 L19 L24 0.00257126
K19_25 L19 L25 0.00372906
K19_26 L19 L26 0.00974585
K19_27 L19 L27 0.00912683
K19_28 L19 L28 0.0045246
K19_29 L19 L29 0.000808
K19_30 L19 L30 0.00227908
K19_31 L19 L31 -9.79653e-05
K19_32 L19 L32 0.0029366
K19_33 L19 L33 0.00475041
K19_34 L19 L34 0.00517634
K19_35 L19 L35 -0.00148153
K19_36 L19 L36 -0.00122744
K19_37 L19 L37 -0.0173051
K19_38 L19 L38 -0.0204891
K20_21 L20 L21 0.0207806
K20_22 L20 L22 0.0176484
K20_23 L20 L23 0.0161682
K20_24 L20 L24 0.00806301
K20_25 L20 L25 0.00676598
K20_26 L20 L26 0.0146033
K20_27 L20 L27 0.0144233
K20_28 L20 L28 0.0132736
K20_29 L20 L29 0.00831361
K20_30 L20 L30 0.00405193
K20_31 L20 L31 -0.0001546
K20_32 L20 L32 0.00103468
K20_33 L20 L33 0.000881108
K20_34 L20 L34 0.000608967
K20_35 L20 L35 -0.00670866
K20_36 L20 L36 -0.00751246
K20_37 L20 L37 -0.00790119
K20_38 L20 L38 -0.0248609
K21_22 L21 L22 0.0326068
K21_23 L21 L23 0.0330523
K21_24 L21 L24 0.0318239
K21_25 L21 L25 0.022967
K21_26 L21 L26 0.0233753
K21_27 L21 L27 0.023351
K21_28 L21 L28 0.0235789
K21_29 L21 L29 0.022359
K21_30 L21 L30 0.0162794
K21_31 L21 L31 -0.00206608
K21_32 L21 L32 -0.00311589
K21_33 L21 L33 -0.00394351
K21_34 L21 L34 -0.00422229
K21_35 L21 L35 -0.0194493
K21_36 L21 L36 -0.0213673
K21_37 L21 L37 -0.0232699
K21_38 L21 L38 -0.024294
K22_23 L22 L23 0.952476
K22_24 L22 L24 0.901892
K22_25 L22 L25 0.849052
K22_26 L22 L26 0.358294
K22_27 L22 L27 0.360083
K22_28 L22 L28 0.35899
K22_29 L22 L29 0.352807
K22_30 L22 L30 0.344651
K22_31 L22 L31 0.00569502
K22_32 L22 L32 0.0162757
K22_33 L22 L33 0.0245001
K22_34 L22 L34 0.0301643
K22_35 L22 L35 0.0419622
K22_36 L22 L36 0.0170068
K22_37 L22 L37 -0.0167204
K22_38 L22 L38 -0.0535464
K23_24 L23 L24 0.946845
K23_25 L23 L25 0.89118
K23_26 L23 L26 0.350553
K23_27 L23 L27 0.352442
K23_28 L23 L28 0.371318
K23_29 L23 L29 0.370002
K23_30 L23 L30 0.361345
K23_31 L23 L31 0.00509932
K23_32 L23 L32 0.0134607
K23_33 L23 L33 0.0190127
K23_34 L23 L34 0.0222155
K23_35 L23 L35 0.0227536
K23_36 L23 L36 0.0172637
K23_37 L23 L37 -0.0110545
K23_38 L23 L38 -0.0482922
K24_25 L24 L25 0.941258
K24_26 L24 L26 0.342819
K24_27 L24 L27 0.344648
K24_28 L24 L28 0.363055
K24_29 L24 L29 0.384115
K24_30 L24 L30 0.380831
K24_31 L24 L31 0.00385007
K24_32 L24 L32 0.00871862
K24_33 L24 L33 0.0113775
K24_34 L24 L34 0.0129197
K24_35 L24 L35 0.00433745
K24_36 L24 L36 0.00149264
K24_37 L24 L37 -0.00595116
K24_38 L24 L38 -0.0374303
K25_26 L25 L26 0.333636
K25_27 L25 L27 0.335439
K25_28 L25 L28 0.353312
K25_29 L25 L29 0.373731
K25_30 L25 L30 0.395737
K25_31 L25 L31 0.00161165
K25_32 L25 L32 0.00319416
K25_33 L25 L33 0.00405255
K25_34 L25 L34 0.00479066
K25_35 L25 L35 -0.00998467
K25_36 L25 L36 -0.0126845
K25_37 L25 L37 -0.0167351
K25_38 L25 L38 -0.024411
K26_27 L26 L27 0.994256
K26_28 L26 L28 0.940864
K26_29 L26 L29 0.884146
K26_30 L26 L30 0.823685
K26_31 L26 L31 0.00511637
K26_32 L26 L32 0.0153032
K26_33 L26 L33 0.0239183
K26_34 L26 L34 0.0305863
K26_35 L26 L35 0.0316251
K26_36 L26 L36 0.0072322
K26_37 L26 L37 -0.0208813
K26_38 L26 L38 -0.0493033
K27_28 L27 L28 0.947016
K27_29 L27 L29 0.889901
K27_30 L27 L30 0.829076
K27_31 L27 L31 0.00485313
K27_32 L27 L32 0.0145906
K27_33 L27 L33 0.0226228
K27_34 L27 L34 0.0285267
K27_35 L27 L35 0.0300335
K27_36 L27 L36 0.00749405
K27_37 L27 L37 -0.0202874
K27_38 L27 L38 -0.0486449
K28_29 L28 L29 0.940658
K28_30 L28 L30 0.876272
K28_31 L28 L31 0.00417137
K28_32 L28 L32 0.0120387
K28_33 L28 L33 0.0177961
K28_34 L28 L34 0.0214055
K28_35 L28 L35 0.0177665
K28_36 L28 L36 0.00849548
K28_37 L28 L37 -0.016284
K28_38 L28 L38 -0.0448618
K29_30 L29 L30 0.932414
K29_31 L29 L31 0.00301464
K29_32 L29 L32 0.00778826
K29_33 L29 L33 0.0107664
K29_34 L29 L34 0.0124849
K29_35 L29 L35 0.00323707
K29_36 L29 L36 0.000105854
K29_37 L29 L37 -0.0104408
K29_38 L29 L38 -0.0357587
K30_31 L30 L31 0.000943055
K30_32 L30 L32 0.00234105
K30_33 L30 L33 0.00315535
K30_34 L30 L34 0.00374111
K30_35 L30 L35 -0.00858045
K30_36 L30 L36 -0.0105618
K30_37 L30 L37 -0.0140154
K30_38 L30 L38 -0.0229545
K31_32 L31 L32 0.467762
K31_33 L31 L33 0.412116
K31_34 L31 L34 0.376285
K31_35 L31 L35 0.316157
K31_36 L31 L36 0.329516
K31_37 L31 L37 0.339538
K31_38 L31 L38 0.340321
K32_33 L32 L33 0.589555
K32_34 L32 L34 0.532103
K32_35 L32 L35 0.337922
K32_36 L32 L36 0.346754
K32_37 L32 L37 0.347235
K32_38 L32 L38 0.33819
K33_34 L33 L34 0.666036
K33_35 L33 L35 0.348101
K33_36 L33 L36 0.349459
K33_37 L33 L37 0.341223
K33_38 L33 L38 0.32785
K34_35 L34 L35 0.347685
K34_36 L34 L36 0.340925
K34_37 L34 L37 0.328216
K34_38 L34 L38 0.313252
K35_36 L35 L36 0.94488
K35_37 L35 L37 0.886734
K35_38 L35 L38 0.825111
K36_37 L36 L37 0.940016
K36_38 L36 L38 0.876367
K37_38 L37 L38 0.935167
.ends Quadraat_series
.ends Quadraat
