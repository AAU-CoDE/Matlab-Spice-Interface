* BEGIN ANSOFT HEADER
* node 1    DC+:D1K
* node 2    DC+:D2K
* node 3    DC+:D3K
* node 4    DC+:D4K
* node 5    DC-:DC-GS-short-b
* node 6    DC-:Q1BW
* node 7    DC-:Q1S
* node 8    DC-:Q2BW
* node 9    DC-:Q2S
* node 10   DC-:Q3BW
* node 11   DC-:Q3S
* node 12   DC-:Q4BW
* node 13   DC-:Q4S
* node 14   DC-:RS1b
* node 15   DC-:RS2b
* node 16   DC-:RS3b
* node 17   DC-:RS4b
* node 18   G1:Q1G
* node 19   G2:Q2G
* node 20   G3:Q3G
* node 21   G4:Q4G
* node 22   GG:RG1a
* node 23   GG:RG2a
* node 24   GG:RG3a
* node 25   GG:RG4a
* node 26   GS:DC-GS-short-a
* node 27   GS:RS1a
* node 28   GS:RS2a
* node 29   GS:RS3a
* node 30   GS:RS4a
* node 31   OUT:D1A
* node 32   OUT:D2A
* node 33   OUT:D3A
* node 34   OUT:D4A
* node 35   OUT:Q1D
* node 36   OUT:Q2D
* node 37   OUT:Q3D
* node 38   OUT:Q4D
* node 39   DC+:DC+terminal
* node 40   DC-:DC-terminal
* node 41   G1:RG1b
* node 42   G2:RG2b
* node 43   G3:RG3b
* node 44   G4:RG4b
* node 45   GG:G-terminal
* node 46   GS:S-terminal
* node 47   OUT:OUT-terminal
*  Project: Quadraat 0004 [4.0 4.0 4.0 4.0]
*   Design: Q3DDesign1
*   Format: Ansys Nexxim
*   Topckt: Quadraat_0004__4_0_4_0_4_0_4
*  Creator: Ansys Electronics Desktop 2022.1.0
*     Date: Wed Nov 30 15:52:13 2022
* END ANSOFT HEADER

.subckt Quadraat 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17
+ 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42 43
+ 44 45 46 47
XZhalf1 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27
+ 28 29 30 31 32 33 34 35 36 37 38 77 78 79 80 81 82 83 84 85 86 87 88 89 90 91
+ 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106 107 108 109 110 111 112
+ 113 114 Quadraat_0004__4_0_4_0_4_0_4_half
XY1 77 78 79 80 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101
+ 102 103 104 105 106 107 108 109 110 111 112 113 114
+ Quadraat_0004__4_0_4_0_4_0_4_parlel
XZhalf2 77 78 79 80 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 39 39 39 39 40 40 40
+ 40 40 40 40 40 40 40 40 40 40 41 42 43 44 45 45 45 45 46 46 46 46 46 47 47 47
+ 47 47 47 47 47 Quadraat_0004__4_0_4_0_4_0_4_half

.subckt Quadraat_0004__4_0_4_0_4_0_4_half 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16
+ 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42
+ 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62 63 64 65 66 67 68
+ 69 70 71 72 73 74 75 76
V1 1 77 dc 0.0
V2 2 78 dc 0.0
V3 3 79 dc 0.0
V4 4 80 dc 0.0
V5 5 81 dc 0.0
V6 6 82 dc 0.0
V7 7 83 dc 0.0
V8 8 84 dc 0.0
V9 9 85 dc 0.0
V10 10 86 dc 0.0
V11 11 87 dc 0.0
V12 12 88 dc 0.0
V13 13 89 dc 0.0
V14 14 90 dc 0.0
V15 15 91 dc 0.0
V16 16 92 dc 0.0
V17 17 93 dc 0.0
V18 18 94 dc 0.0
V19 19 95 dc 0.0
V20 20 96 dc 0.0
V21 21 97 dc 0.0
V22 22 98 dc 0.0
V23 23 99 dc 0.0
V24 24 100 dc 0.0
V25 25 101 dc 0.0
V26 26 102 dc 0.0
V27 27 103 dc 0.0
V28 28 104 dc 0.0
V29 29 105 dc 0.0
V30 30 106 dc 0.0
V31 31 107 dc 0.0
V32 32 108 dc 0.0
V33 33 109 dc 0.0
V34 34 110 dc 0.0
V35 35 111 dc 0.0
V36 36 112 dc 0.0
V37 37 113 dc 0.0
V38 38 114 dc 0.0
R1 77 115 0.00051090800525
R2 78 116 0.000487621597364
R3 79 117 0.000464125221666
R4 80 118 0.000440757961714
R5 81 119 0.000802359878137
R6 82 120 0.000496997612507
R7 83 121 0.0012954071055
R8 84 122 0.000540709589976
R9 85 123 0.00134184790636
R10 86 124 0.000582354317808
R11 87 125 0.00137837008649
R12 88 126 0.00062141584397
R13 89 127 0.0014210443183
R14 90 128 0.00328703345681
R15 91 129 0.00333603995144
R16 92 130 0.00336505616913
R17 93 131 0.00341484227782
R18 94 132 0.00182942294249
R19 95 133 0.00182526969824
R20 96 134 0.00182780123238
R21 97 135 0.00183247816993
R22 98 136 0.0025146969477
R23 99 137 0.00231254669589
R24 100 138 0.00211077600234
R25 101 139 0.00190889671467
R26 102 140 0.00270896308861
R27 103 141 0.00232892322555
R28 104 142 0.00212924727201
R29 105 143 0.00192855472492
R30 106 144 0.00172822643075
R31 107 145 0.00157772338845
R32 108 146 0.00163736558864
R33 109 147 0.00170007496605
R34 110 148 0.00175960912344
R35 111 149 0.000929601117745
R36 112 150 0.000907180444568
R37 113 151 0.000884671709108
R38 114 152 0.00086282768782
F1_2 115 77 V2 0.954075
F1_3 115 77 V3 0.908105
F1_4 115 77 V4 0.862443
F2_1 116 78 V1 0.999637
F2_3 116 78 V3 0.951471
F2_4 116 78 V4 0.903629
F3_1 117 79 V1 0.999639
F3_2 117 79 V2 0.99964
F3_4 117 79 V4 0.949376
F4_1 118 80 V1 0.999708
F4_2 118 80 V2 0.999708
F4_3 118 80 V3 0.999708
F5_6 119 81 V6 0.512053
F5_7 119 81 V7 0.512054
F5_8 119 81 V8 0.512048
F5_9 119 81 V9 0.512048
F5_10 119 81 V10 0.512048
F5_11 119 81 V11 0.512048
F5_12 119 81 V12 0.512048
F5_13 119 81 V13 0.512048
F5_14 119 81 V14 0.512054
F5_15 119 81 V15 0.512048
F5_16 119 81 V16 0.512048
F5_17 119 81 V17 0.512048
F6_5 120 82 V5 0.826666
F6_7 120 82 V7 0.996216
F6_8 120 82 V8 0.979534
F6_9 120 82 V9 0.979538
F6_10 120 82 V10 0.979372
F6_11 120 82 V11 0.979372
F6_12 120 82 V12 0.97937
F6_13 120 82 V13 0.97937
F6_14 120 82 V14 0.996216
F6_15 120 82 V15 0.979538
F6_16 120 82 V16 0.979372
F6_17 120 82 V17 0.97937
F7_5 121 83 V5 0.31716
F7_6 121 83 V6 0.38221
F7_8 121 83 V8 0.375828
F7_9 121 83 V9 0.375829
F7_10 121 83 V10 0.375764
F7_11 121 83 V11 0.375764
F7_12 121 83 V12 0.375763
F7_13 121 83 V13 0.375763
F7_14 121 83 V14 1.00004
F7_15 121 83 V15 0.375829
F7_16 121 83 V16 0.375764
F7_17 121 83 V17 0.375763
F8_5 122 84 V5 0.75983
F8_6 122 84 V6 0.900347
F8_7 122 84 V7 0.900391
F8_9 122 84 V9 0.993829
F8_10 122 84 V10 0.976733
F8_11 122 84 V11 0.976736
F8_12 122 84 V12 0.976571
F8_13 122 84 V13 0.976572
F8_14 122 84 V14 0.900392
F8_15 122 84 V15 0.993829
F8_16 122 84 V16 0.976736
F8_17 122 84 V17 0.976572
F9_5 123 85 V5 0.30618
F9_6 123 85 V6 0.362804
F9_7 123 85 V7 0.362822
F9_8 123 85 V8 0.400472
F9_10 123 85 V10 0.3936
F9_11 123 85 V11 0.393602
F9_12 123 85 V12 0.393534
F9_13 123 85 V13 0.393534
F9_14 123 85 V14 0.362822
F9_15 123 85 V15 1
F9_16 123 85 V16 0.393602
F9_17 123 85 V17 0.393534
F10_5 124 86 V5 0.705493
F10_6 124 86 V6 0.835824
F10_7 124 86 V7 0.835861
F10_8 124 86 V8 0.906886
F10_9 124 86 V9 0.906925
F10_11 124 86 V11 0.993568
F10_12 124 86 V12 0.977369
F10_13 124 86 V13 0.977374
F10_14 124 86 V14 0.835861
F10_15 124 86 V15 0.906925
F10_16 124 86 V16 0.993568
F10_17 124 86 V17 0.977374
F11_5 125 87 V5 0.298067
F11_6 125 87 V6 0.353131
F11_7 125 87 V7 0.353147
F11_8 125 87 V8 0.383156
F11_9 125 87 V9 0.383172
F11_10 125 87 V10 0.419778
F11_12 125 87 V12 0.412944
F11_13 125 87 V13 0.412946
F11_14 125 87 V14 0.353147
F11_15 125 87 V15 0.383172
F11_16 125 87 V16 1
F11_17 125 87 V17 0.412946
F12_5 126 88 V5 0.661147
F12_6 126 88 V6 0.783283
F12_7 126 88 V7 0.783318
F12_8 126 88 V8 0.849739
F12_9 126 88 V9 0.849773
F12_10 126 88 V10 0.915933
F12_11 126 88 V11 0.915957
F12_13 126 88 V13 0.998017
F12_14 126 88 V14 0.783318
F12_15 126 88 V15 0.849773
F12_16 126 88 V16 0.915957
F12_17 126 88 V17 0.998017
F13_5 127 89 V5 0.289116
F13_6 127 89 V6 0.342526
F13_7 127 89 V7 0.342541
F13_8 127 89 V8 0.371587
F13_9 127 89 V9 0.371602
F13_10 127 89 V10 0.400535
F13_11 127 89 V11 0.400545
F13_12 127 89 V12 0.436428
F13_14 127 89 V14 0.342541
F13_15 127 89 V15 0.371602
F13_16 127 89 V16 0.400545
F13_17 127 89 V17 0.999999
F14_5 128 90 V5 0.124991
F14_6 128 90 V6 0.150627
F14_7 128 90 V7 0.394111
F14_8 128 90 V8 0.148112
F14_9 128 90 V9 0.148113
F14_10 128 90 V10 0.148087
F14_11 128 90 V11 0.148087
F14_12 128 90 V12 0.148087
F14_13 128 90 V13 0.148087
F14_15 128 90 V15 0.148113
F14_16 128 90 V16 0.148087
F14_17 128 90 V17 0.148087
F15_5 129 91 V5 0.123154
F15_6 129 91 V6 0.14593
F15_7 129 91 V7 0.145937
F15_8 129 91 V8 0.161081
F15_9 129 91 V9 0.402228
F15_10 129 91 V10 0.158317
F15_11 129 91 V11 0.158317
F15_12 129 91 V12 0.15829
F15_13 129 91 V13 0.15829
F15_14 129 91 V14 0.145937
F15_16 129 91 V16 0.158317
F15_17 129 91 V17 0.15829
F16_5 130 92 V5 0.122092
F16_6 130 92 V6 0.144647
F16_7 130 92 V7 0.144654
F16_8 130 92 V8 0.156946
F16_9 130 92 V9 0.156952
F16_10 130 92 V10 0.171946
F16_11 130 92 V11 0.409613
F16_12 130 92 V12 0.169147
F16_13 130 92 V13 0.169148
F16_14 130 92 V14 0.144654
F16_15 130 92 V15 0.156952
F16_17 130 92 V17 0.169148
F17_5 131 93 V5 0.120312
F17_6 131 93 V6 0.142538
F17_7 131 93 V7 0.142544
F17_8 131 93 V8 0.154631
F17_9 131 93 V9 0.154637
F17_10 131 93 V10 0.166678
F17_11 131 93 V11 0.166682
F17_12 131 93 V12 0.181614
F17_13 131 93 V13 0.416137
F17_14 131 93 V14 0.142544
F17_15 131 93 V15 0.154637
F17_16 131 93 V16 0.166682
F22_23 136 98 V23 0.919593
F22_24 136 98 V24 0.839358
F22_25 136 98 V25 0.759075
F23_22 137 99 V22 0.999979
F23_24 137 99 V24 0.91273
F23_25 137 99 V25 0.82543
F24_22 138 100 V22 0.999979
F24_23 138 100 V23 0.999979
F24_25 138 100 V25 0.904333
F25_22 139 101 V22 0.999973
F25_23 139 101 V23 0.999973
F25_24 139 101 V24 0.999973
F26_27 140 102 V27 0.859685
F26_28 140 102 V28 0.785988
F26_29 140 102 V29 0.711899
F26_30 140 102 V30 0.637952
F27_26 141 103 V26 0.999971
F27_28 141 103 V28 0.914248
F27_29 141 103 V29 0.828069
F27_30 141 103 V30 0.742055
F28_26 142 104 V26 0.999984
F28_27 142 104 V27 0.999984
F28_29 142 104 V29 0.905724
F28_30 142 104 V30 0.811643
F29_26 143 105 V26 0.999977
F29_27 143 105 V27 0.999977
F29_28 143 105 V28 0.999977
F29_30 143 105 V30 0.896106
F30_26 144 106 V26 0.999978
F30_27 144 106 V27 0.999978
F30_28 144 106 V28 0.999978
F30_29 144 106 V29 0.999978
F31_32 145 107 V32 0.493496
F31_33 145 107 V33 0.493503
F31_34 145 107 V34 0.493503
F31_35 145 107 V35 0.464197
F31_36 145 107 V36 0.464197
F31_37 145 107 V37 0.464197
F31_38 145 107 V38 0.464197
F32_31 146 108 V31 0.47552
F32_33 146 108 V33 0.513057
F32_34 146 108 V34 0.513056
F32_35 146 108 V35 0.447306
F32_36 146 108 V36 0.447306
F32_37 146 108 V37 0.447306
F32_38 146 108 V38 0.447306
F33_31 147 109 V31 0.457986
F33_32 147 109 V32 0.494132
F33_34 147 109 V34 0.530259
F33_35 147 109 V35 0.430807
F33_36 147 109 V36 0.430807
F33_37 147 109 V37 0.430807
F33_38 147 109 V38 0.430806
F34_31 148 110 V31 0.442491
F34_32 148 110 V32 0.477413
F34_33 148 110 V33 0.512318
F34_35 148 110 V35 0.416231
F34_36 148 110 V36 0.416231
F34_37 148 110 V37 0.416231
F34_38 148 110 V38 0.416231
F35_31 149 111 V31 0.787838
F35_32 149 111 V32 0.787868
F35_33 149 111 V33 0.787868
F35_34 149 111 V34 0.787868
F35_36 149 111 V36 0.975111
F35_37 149 111 V37 0.950902
F35_38 149 111 V38 0.927115
F36_31 150 112 V31 0.807309
F36_32 150 112 V32 0.80734
F36_33 150 112 V33 0.80734
F36_34 150 112 V34 0.80734
F36_35 150 112 V35 0.99921
F36_37 150 112 V37 0.974406
F36_38 150 112 V38 0.950028
F37_31 151 113 V31 0.827849
F37_32 151 113 V32 0.827881
F37_33 151 113 V33 0.827882
F37_34 151 113 V34 0.827882
F37_35 151 113 V35 0.999195
F37_36 151 113 V36 0.999198
F37_38 151 113 V38 0.974203
F38_31 152 114 V31 0.848808
F38_32 152 114 V32 0.848841
F38_33 152 114 V33 0.848841
F38_34 152 114 V34 0.848841
F38_35 152 114 V35 0.998864
F38_36 152 114 V36 0.998864
F38_37 152 114 V37 0.998867
L1 115 39 4.91154680987e-09
L2 116 40 4.57697651557e-09
L3 117 41 4.22784815784e-09
L4 118 42 3.8370363576e-09
L5 119 43 3.76508702107e-09
L6 120 44 4.41190769607e-09
L7 121 45 5.35487424543e-09
L8 122 46 5.05811970061e-09
L9 123 47 6.05992206174e-09
L10 124 48 5.66670328607e-09
L11 125 49 6.69390947072e-09
L12 126 50 6.30375567286e-09
L13 127 51 7.34249491902e-09
L14 128 52 7.26947181218e-09
L15 129 53 8.03154867793e-09
L16 130 54 8.68325922631e-09
L17 131 55 9.33366268216e-09
L18 132 56 1.80713680406e-09
L19 133 57 1.81432100611e-09
L20 134 58 1.81488117957e-09
L21 135 59 1.82467587804e-09
L22 136 60 7.78541235511e-09
L23 137 61 6.99144742317e-09
L24 138 62 6.18817045926e-09
L25 139 63 5.39367081581e-09
L26 140 64 8.65562703106e-09
L27 141 65 8.27724216315e-09
L28 142 66 7.40492457149e-09
L29 143 67 6.52754978448e-09
L30 144 68 5.63056302677e-09
L31 145 69 5.97335049799e-09
L32 146 70 6.57569021799e-09
L33 147 71 7.27974699819e-09
L34 148 72 8.04182617335e-09
L35 149 73 7.34886754509e-09
L36 150 74 7.09809709956e-09
L37 151 75 6.9244110772e-09
L38 152 76 6.84828363478e-09
K1_2 L1 L2 0.97011
K1_3 L1 L3 0.937523
K1_4 L1 L4 0.902755
K1_5 L1 L5 0.138467
K1_6 L1 L6 0.135215
K1_7 L1 L7 0.129078
K1_8 L1 L8 0.158757
K1_9 L1 L9 0.144933
K1_10 L1 L10 0.173807
K1_11 L1 L11 0.155788
K1_12 L1 L12 0.17987
K1_13 L1 L13 0.160785
K1_14 L1 L14 0.11201
K1_15 L1 L15 0.125229
K1_16 L1 L16 0.134984
K1_17 L1 L17 0.140033
K1_18 L1 L18 -0.00735397
K1_19 L1 L19 -0.00358714
K1_20 L1 L20 -0.000670389
K1_21 L1 L21 0.00142309
K1_22 L1 L22 0.00296039
K1_23 L1 L23 0.0129222
K1_24 L1 L24 0.0226728
K1_25 L1 L25 0.0311221
K1_26 L1 L26 -0.0120557
K1_27 L1 L27 -0.004788
K1_28 L1 L28 0.00433801
K1_29 L1 L29 0.0134931
K1_30 L1 L30 0.0217944
K1_31 L1 L31 0.0435892
K1_32 L1 L32 0.00702323
K1_33 L1 L33 -0.0327882
K1_34 L1 L34 -0.0750596
K1_35 L1 L35 -0.019653
K1_36 L1 L36 -0.00485904
K1_37 L1 L37 0.00770244
K1_38 L1 L38 0.0167675
K2_3 L2 L3 0.967818
K2_4 L2 L4 0.932224
K2_5 L2 L5 0.139486
K2_6 L2 L6 0.138829
K2_7 L2 L7 0.130907
K2_8 L2 L8 0.160138
K2_9 L2 L9 0.144787
K2_10 L2 L10 0.169098
K2_11 L2 L11 0.151685
K2_12 L2 L12 0.169079
K2_13 L2 L13 0.152777
K2_14 L2 L14 0.113096
K2_15 L2 L15 0.124811
K2_16 L2 L16 0.131552
K2_17 L2 L17 0.133609
K2_18 L2 L18 -0.00616532
K2_19 L2 L19 -0.00240899
K2_20 L2 L20 -0.000165702
K2_21 L2 L21 0.000887409
K2_22 L2 L22 0.00698612
K2_23 L2 L23 0.0160745
K2_24 L2 L24 0.0242997
K2_25 L2 L25 0.0311707
K2_26 L2 L26 -0.00739014
K2_27 L2 L27 -0.000200199
K2_28 L2 L28 0.00830139
K2_29 L2 L29 0.0162582
K2_30 L2 L30 0.0231841
K2_31 L2 L31 0.0400193
K2_32 L2 L32 0.0283485
K2_33 L2 L33 -0.00883162
K2_34 L2 L34 -0.0530544
K2_35 L2 L35 -0.00936975
K2_36 L2 L36 0.00423278
K2_37 L2 L37 0.0142906
K2_38 L2 L38 0.0206452
K3_4 L3 L4 0.964758
K3_5 L3 L5 0.139109
K3_6 L3 L6 0.14205
K3_7 L3 L7 0.131674
K3_8 L3 L8 0.157317
K3_9 L3 L9 0.141589
K3_10 L3 L10 0.159307
K3_11 L3 L11 0.14407
K3_12 L3 L12 0.156636
K3_13 L3 L13 0.14295
K3_14 L3 L14 0.113082
K3_15 L3 L15 0.121902
K3_16 L3 L16 0.125274
K3_17 L3 L17 0.125517
K3_18 L3 L18 -0.00445803
K3_19 L3 L19 -0.00135488
K3_20 L3 L20 -0.000103115
K3_21 L3 L21 0.000307252
K3_22 L3 L22 0.0116357
K3_23 L3 L23 0.0193714
K3_24 L3 L24 0.0259216
K3_25 L3 L25 0.0315319
K3_26 L3 L26 -0.00202986
K3_27 L3 L27 0.0049079
K3_28 L3 L28 0.0123864
K3_29 L3 L29 0.0189172
K3_30 L3 L30 0.02462
K3_31 L3 L31 0.0413298
K3_32 L3 L32 0.0348291
K3_33 L3 L33 0.0214676
K3_34 L3 L34 -0.0207719
K3_35 L3 L35 0.00685944
K3_36 L3 L36 0.0182374
K3_37 L3 L37 0.0254885
K3_38 L3 L38 0.0299641
K4_5 L4 L5 0.13667
K4_6 L4 L6 0.14188
K4_7 L4 L7 0.129741
K4_8 L4 L8 0.148846
K4_9 L4 L9 0.134632
K4_10 L4 L10 0.147355
K4_11 L4 L11 0.134402
K4_12 L4 L12 0.143829
K4_13 L4 L13 0.132221
K4_14 L4 L14 0.110793
K4_15 L4 L15 0.115987
K4_16 L4 L16 0.117202
K4_17 L4 L17 0.116442
K4_18 L4 L18 -0.00263785
K4_19 L4 L19 -0.000745159
K4_20 L4 L20 -0.000193434
K4_21 L4 L21 -7.18044e-05
K4_22 L4 L22 0.0162586
K4_23 L4 L23 0.0224661
K4_24 L4 L24 0.0276812
K4_25 L4 L25 0.0324324
K4_26 L4 L26 0.00353434
K4_27 L4 L27 0.010036
K4_28 L4 L28 0.0162642
K4_29 L4 L29 0.0215397
K4_30 L4 L30 0.0263492
K4_31 L4 L31 0.0446014
K4_32 L4 L32 0.0386795
K4_33 L4 L33 0.0304013
K4_34 L4 L34 0.0118659
K4_35 L4 L35 0.0213463
K4_36 L4 L36 0.029879
K4_37 L4 L37 0.0350655
K4_38 L4 L38 0.0383827
K5_6 L5 L6 0.802868
K5_7 L5 L7 0.737008
K5_8 L5 L8 0.76627
K5_9 L5 L9 0.704635
K5_10 L5 L10 0.72982
K5_11 L5 L11 0.674496
K5_12 L5 L12 0.695347
K5_13 L5 L13 0.646337
K5_14 L5 L14 0.637558
K5_15 L5 L15 0.614507
K5_16 L5 L16 0.593525
K5_17 L5 L17 0.574008
K5_18 L5 L18 -0.0134941
K5_19 L5 L19 -0.00516006
K5_20 L5 L20 -0.00297224
K5_21 L5 L21 -0.00249815
K5_22 L5 L22 0.0250674
K5_23 L5 L23 0.0284785
K5_24 L5 L24 0.0315557
K5_25 L5 L25 0.0352157
K5_26 L5 L26 -0.00167004
K5_27 L5 L27 0.0171233
K5_28 L5 L28 0.0219669
K5_29 L5 L29 0.0251345
K5_30 L5 L30 0.0286871
K5_31 L5 L31 0.0347476
K5_32 L5 L32 0.0278822
K5_33 L5 L33 0.0190738
K5_34 L5 L34 0.00693786
K5_35 L5 L35 0.0299281
K5_36 L5 L36 0.0388188
K5_37 L5 L37 0.0422487
K5_38 L5 L38 0.044379
K6_7 L6 L7 0.893921
K6_8 L6 L8 0.933061
K6_9 L6 L9 0.845815
K6_10 L6 L10 0.883565
K6_11 L6 L11 0.809339
K6_12 L6 L12 0.840549
K6_13 L6 L13 0.776244
K6_14 L6 L14 0.751921
K6_15 L6 L15 0.728875
K6_16 L6 L16 0.707775
K6_17 L6 L17 0.686492
K6_18 L6 L18 0.00931858
K6_19 L6 L19 0.00449629
K6_20 L6 L20 0.00247101
K6_21 L6 L21 0.00179776
K6_22 L6 L22 0.0115005
K6_23 L6 L23 0.0265037
K6_24 L6 L24 0.0347877
K6_25 L6 L25 0.0409586
K6_26 L6 L26 -0.0222587
K6_27 L6 L27 -0.00342071
K6_28 L6 L28 0.0154916
K6_29 L6 L29 0.0254339
K6_30 L6 L30 0.0321703
K6_31 L6 L31 0.0238038
K6_32 L6 L32 0.0211968
K6_33 L6 L33 0.0174486
K6_34 L6 L34 0.00683349
K6_35 L6 L35 -0.0115721
K6_36 L6 L36 0.00188458
K6_37 L6 L37 0.00721063
K6_38 L6 L38 0.0105668
K7_8 L7 L8 0.834924
K7_9 L7 L9 0.765702
K7_10 L7 L10 0.791311
K7_11 L7 L11 0.72851
K7_12 L7 L12 0.75293
K7_13 L7 L13 0.697705
K7_14 L7 L14 0.847081
K7_15 L7 L15 0.663597
K7_16 L7 L16 0.638998
K7_17 L7 L17 0.618312
K7_18 L7 L18 0.00542808
K7_19 L7 L19 -0.000360743
K7_20 L7 L20 -0.000393246
K7_21 L7 L21 -0.000504655
K7_22 L7 L22 0.0136582
K7_23 L7 L23 0.0249748
K7_24 L7 L24 0.0308536
K7_25 L7 L25 0.0355855
K7_26 L7 L26 -0.0179979
K7_27 L7 L27 9.68748e-05
K7_28 L7 L28 0.0157081
K7_29 L7 L29 0.0230583
K7_30 L7 L30 0.0281529
K7_31 L7 L31 0.027143
K7_32 L7 L32 0.0220886
K7_33 L7 L33 0.0151679
K7_34 L7 L34 0.00313887
K7_35 L7 L35 0.0126681
K7_36 L7 L36 0.0212814
K7_37 L7 L37 0.0248099
K7_38 L7 L38 0.0272588
K8_9 L8 L9 0.90728
K8_10 L8 L10 0.940796
K8_11 L8 L11 0.861872
K8_12 L8 L12 0.893835
K8_13 L8 L13 0.82592
K8_14 L8 L14 0.704041
K8_15 L8 L15 0.780943
K8_16 L8 L16 0.752998
K8_17 L8 L17 0.730356
K8_18 L8 L18 0.00181339
K8_19 L8 L19 0.00331167
K8_20 L8 L20 0.00251605
K8_21 L8 L21 0.00144903
K8_22 L8 L22 -0.00378318
K8_23 L8 L23 0.0193938
K8_24 L8 L24 0.0313408
K8_25 L8 L25 0.0387085
K8_26 L8 L26 -0.0385203
K8_27 L8 L27 -0.0187535
K8_28 L8 L28 0.00590477
K8_29 L8 L29 0.0202402
K8_30 L8 L30 0.0287199
K8_31 L8 L31 0.0256003
K8_32 L8 L32 0.0190171
K8_33 L8 L33 0.00465756
K8_34 L8 L34 -0.0194742
K8_35 L8 L35 -0.0301775
K8_36 L8 L36 0.00423271
K8_37 L8 L37 0.0138505
K8_38 L8 L38 0.017841
K9_10 L9 L10 0.853991
K9_11 L9 L11 0.790056
K9_12 L9 L12 0.812024
K9_13 L9 L13 0.75367
K9_14 L9 L14 0.64899
K9_15 L9 L15 0.863596
K9_16 L9 L16 0.693449
K9_17 L9 L17 0.668208
K9_18 L9 L18 -0.00500737
K9_19 L9 L19 0.00112147
K9_20 L9 L20 -0.00178058
K9_21 L9 L21 -0.00148576
K9_22 L9 L22 -0.00308557
K9_23 L9 L23 0.0189375
K9_24 L9 L24 0.0281828
K9_25 L9 L25 0.0338218
K9_26 L9 L26 -0.0357089
K9_27 L9 L27 -0.0168563
K9_28 L9 L28 0.00642302
K9_29 L9 L29 0.0187116
K9_30 L9 L30 0.0253293
K9_31 L9 L31 0.0281474
K9_32 L9 L32 0.0193608
K9_33 L9 L33 0.00524204
K9_34 L9 L34 -0.0152175
K9_35 L9 L35 -0.0072628
K9_36 L9 L36 0.0278965
K9_37 L9 L37 0.0334934
K9_38 L9 L38 0.0361968
K10_11 L10 L11 0.916422
K10_12 L10 L12 0.945366
K10_13 L10 L13 0.873387
K10_14 L10 L14 0.668194
K10_15 L10 L15 0.736131
K10_16 L10 L16 0.799395
K10_17 L10 L17 0.771422
K10_18 L10 L18 -0.00143217
K10_19 L10 L19 -0.00257001
K10_20 L10 L20 0.00177958
K10_21 L10 L21 0.00172442
K10_22 L10 L22 -0.0204829
K10_23 L10 L23 0.00571703
K10_24 L10 L24 0.026322
K10_25 L10 L25 0.0376555
K10_26 L10 L26 -0.0542403
K10_27 L10 L27 -0.035022
K10_28 L10 L28 -0.00875231
K10_29 L10 L29 0.0118846
K10_30 L10 L30 0.025017
K10_31 L10 L31 0.0289503
K10_32 L10 L32 0.0102255
K10_33 L10 L33 -0.0162133
K10_34 L10 L34 -0.0432408
K10_35 L10 L35 -0.0433587
K10_36 L10 L36 -0.00667074
K10_37 L10 L37 0.0232225
K10_38 L10 L38 0.0315622
K11_12 L11 L12 0.866917
K11_13 L11 L13 0.808297
K11_14 L11 L14 0.616963
K11_15 L11 L15 0.683644
K11_16 L11 L16 0.874527
K11_17 L11 L17 0.717076
K11_18 L11 L18 -0.00472287
K11_19 L11 L19 -0.00844004
K11_20 L11 L20 -0.000358855
K11_21 L11 L21 -0.00304894
K11_22 L11 L22 -0.0218436
K11_23 L11 L23 0.0033836
K11_24 L11 L24 0.0236513
K11_25 L11 L25 0.032953
K11_26 L11 L26 -0.0531512
K11_27 L11 L27 -0.0350218
K11_28 L11 L28 -0.0100606
K11_29 L11 L29 0.0101749
K11_30 L11 L30 0.0219453
K11_31 L11 L31 0.0297449
K11_32 L11 L32 0.0127479
K11_33 L11 L33 -0.00928526
K11_34 L11 L34 -0.0325464
K11_35 L11 L35 -0.0189644
K11_36 L11 L36 0.0164295
K11_37 L11 L37 0.0478236
K11_38 L11 L38 0.0526827
K12_13 L12 L13 0.923603
K12_14 L12 L14 0.636057
K12_15 L12 L15 0.70067
K12_16 L12 L16 0.757058
K12_17 L12 L17 0.81399
K12_18 L12 L18 -0.00247984
K12_19 L12 L19 -0.00528108
K12_20 L12 L20 -0.00357026
K12_21 L12 L21 0.00183802
K12_22 L12 L22 -0.0326979
K12_23 L12 L23 -0.00678805
K12_24 L12 L24 0.0173857
K12_25 L12 L25 0.0376987
K12_26 L12 L26 -0.0663276
K12_27 L12 L27 -0.0480439
K12_28 L12 L28 -0.0224343
K12_29 L12 L29 0.000294662
K12_30 L12 L30 0.0199321
K12_31 L12 L31 0.026958
K12_32 L12 L32 -0.00327811
K12_33 L12 L33 -0.0320178
K12_34 L12 L34 -0.0584887
K12_35 L12 L35 -0.0449218
K12_36 L12 L36 -0.00940751
K12_37 L12 L37 0.0233255
K12_38 L12 L38 0.0521261
K13_14 L13 L14 0.590628
K13_15 L13 L15 0.651818
K13_16 L13 L16 0.708429
K13_17 L13 L17 0.883972
K13_18 L13 L18 -0.00451542
K13_19 L13 L19 -0.00816631
K13_20 L13 L20 -0.00963635
K13_21 L13 L21 -0.00201804
K13_22 L13 L22 -0.0361952
K13_23 L13 L23 -0.0116246
K13_24 L13 L24 0.0122407
K13_25 L13 L25 0.0330189
K13_26 L13 L26 -0.0671503
K13_27 L13 L27 -0.049983
K13_28 L13 L28 -0.025885
K13_29 L13 L29 -0.00369492
K13_30 L13 L30 0.0162382
K13_31 L13 L31 0.0285025
K13_32 L13 L32 0.00381636
K13_33 L13 L33 -0.0207367
K13_34 L13 L34 -0.0443063
K13_35 L13 L35 -0.0131778
K13_36 L13 L36 0.0209959
K13_37 L13 L37 0.0531713
K13_38 L13 L38 0.0837355
K14_15 L14 L15 0.568965
K14_16 L14 L16 0.542919
K14_17 L14 L17 0.524348
K14_18 L14 L18 -0.118278
K14_19 L14 L19 -0.00778262
K14_20 L14 L20 -0.00277494
K14_21 L14 L21 -0.00194764
K14_22 L14 L22 0.0148047
K14_23 L14 L23 0.0213329
K14_24 L14 L24 0.0251166
K14_25 L14 L25 0.0285934
K14_26 L14 L26 -0.0166701
K14_27 L14 L27 0.00437999
K14_28 L14 L28 0.014657
K14_29 L14 L29 0.0192163
K14_30 L14 L30 0.0228128
K14_31 L14 L31 0.0255695
K14_32 L14 L32 0.0203714
K14_33 L14 L33 0.0134479
K14_34 L14 L34 0.00236172
K14_35 L14 L35 0.0166456
K14_36 L14 L36 0.0259414
K14_37 L14 L37 0.0291274
K14_38 L14 L38 0.0311118
K15_16 L15 L16 0.605638
K15_17 L15 L17 0.57945
K15_18 L15 L18 -0.0207277
K15_19 L15 L19 -0.114207
K15_20 L15 L20 -0.00825047
K15_21 L15 L21 -0.00364044
K15_22 L15 L22 -0.00112094
K15_23 L15 L23 0.0179135
K15_24 L15 L24 0.0232899
K15_25 L15 L25 0.0272329
K15_26 L15 L26 -0.0309986
K15_27 L15 L27 -0.0136181
K15_28 L15 L28 0.00780118
K15_29 L15 L29 0.0163416
K15_30 L15 L30 0.0207232
K15_31 L15 L31 0.0261746
K15_32 L15 L32 0.0180148
K15_33 L15 L33 0.00556236
K15_34 L15 L34 -0.0119688
K15_35 L15 L35 0.00195969
K15_36 L15 L36 0.0293152
K15_37 L15 L37 0.0360302
K15_38 L15 L38 0.0386351
K16_17 L16 L17 0.633831
K16_18 L16 L18 -0.00759925
K16_19 L16 L19 -0.0227544
K16_20 L16 L20 -0.111144
K16_21 L16 L21 -0.00963802
K16_22 L16 L22 -0.0214664
K16_23 L16 L23 0.00169094
K16_24 L16 L24 0.0195878
K16_25 L16 L25 0.0251729
K16_26 L16 L26 -0.0489953
K16_27 L16 L27 -0.0327522
K16_28 L16 L28 -0.0101156
K16_29 L16 L29 0.00920553
K16_30 L16 L30 0.0175105
K16_31 L16 L31 0.0274851
K16_32 L16 L32 0.0127906
K16_33 L16 L33 -0.00599737
K16_34 L16 L34 -0.025934
K16_35 L16 L35 -0.00783958
K16_36 L16 L36 0.0229287
K16_37 L16 L37 0.0474178
K16_38 L16 L38 0.0535397
K17_18 L17 L18 -0.00566872
K17_19 L17 L19 -0.0106063
K17_20 L17 L20 -0.0237289
K17_21 L17 L21 -0.110013
K17_22 L17 L22 -0.042599
K17_23 L17 L23 -0.0208947
K17_24 L17 L24 0.00109149
K17_25 L17 L25 0.0195314
K17_26 L17 L26 -0.066755
K17_27 L17 L27 -0.0514885
K17_28 L17 L28 -0.0301415
K17_29 L17 L29 -0.00973856
K17_30 L17 L30 0.00952242
K17_31 L17 L31 0.0267389
K17_32 L17 L32 0.00588681
K17_33 L17 L33 -0.01513
K17_34 L17 L34 -0.0356196
K17_35 L17 L35 -0.00148229
K17_36 L17 L36 0.0291036
K17_37 L17 L37 0.0573882
K17_38 L17 L38 0.0813941
K18_19 L18 L19 0.0189789
K18_20 L18 L20 0.00506591
K18_21 L18 L21 0.00293585
K18_22 L18 L22 0.000538625
K18_23 L18 L23 0.000338114
K18_24 L18 L24 0.00183892
K18_25 L18 L25 0.00244381
K18_26 L18 L26 0.00767422
K18_27 L18 L27 0.00203503
K18_28 L18 L28 -0.000362067
K18_29 L18 L29 0.00139309
K18_30 L18 L30 0.00226401
K18_31 L18 L31 -0.00381072
K18_32 L18 L32 -0.00160957
K18_33 L18 L33 0.000972051
K18_34 L18 L34 0.00327243
K18_35 L18 L35 -0.00236407
K18_36 L18 L36 -0.0122118
K18_37 L18 L37 -0.0138238
K18_38 L18 L38 -0.0141348
K19_20 L19 L20 0.0186195
K19_21 L19 L21 0.00542665
K19_22 L19 L22 0.00984257
K19_23 L19 L23 0.00314641
K19_24 L19 L24 0.00141918
K19_25 L19 L25 0.00247613
K19_26 L19 L26 0.00975439
K19_27 L19 L27 0.0085533
K19_28 L19 L28 0.00448551
K19_29 L19 L29 0.000775278
K19_30 L19 L30 0.00208752
K19_31 L19 L31 -0.00345883
K19_32 L19 L32 -0.00136433
K19_33 L19 L33 0.000167991
K19_34 L19 L34 0.000822952
K19_35 L19 L35 -0.00422721
K19_36 L19 L36 -0.00427003
K19_37 L19 L37 -0.0142081
K19_38 L19 L38 -0.0159773
K20_21 L20 L21 0.0199989
K20_22 L20 L22 0.0158374
K20_23 L20 L23 0.0144545
K20_24 L20 L24 0.00708284
K20_25 L20 L25 0.00490058
K20_26 L20 L26 0.0139419
K20_27 L20 L27 0.0136421
K20_28 L20 L28 0.0126544
K20_29 L20 L29 0.00803242
K20_30 L20 L30 0.00384406
K20_31 L20 L31 -0.00287238
K20_32 L20 L32 -0.00192338
K20_33 L20 L33 -0.00181886
K20_34 L20 L34 -0.00192366
K20_35 L20 L35 -0.0070212
K20_36 L20 L36 -0.00749316
K20_37 L20 L37 -0.00769647
K20_38 L20 L38 -0.0179153
K21_22 L21 L22 0.0224488
K21_23 L21 L23 0.0225409
K21_24 L21 L24 0.0207906
K21_25 L21 L25 0.0116285
K21_26 L21 L26 0.0213911
K21_27 L21 L27 0.0214421
K21_28 L21 L28 0.0216843
K21_29 L21 L29 0.0204918
K21_30 L21 L30 0.0148484
K21_31 L21 L31 -0.00324792
K21_32 L21 L32 -0.003974
K21_33 L21 L33 -0.0045846
K21_34 L21 L34 -0.00483927
K21_35 L21 L35 -0.0148758
K21_36 L21 L36 -0.0157893
K21_37 L21 L37 -0.016628
K21_38 L21 L38 -0.0170749
K22_23 L22 L23 0.94789
K22_24 L22 L24 0.892708
K22_25 L22 L25 0.833625
K22_26 L22 L26 0.307851
K22_27 L22 L27 0.316528
K22_28 L22 L28 0.313267
K22_29 L22 L29 0.305365
K22_30 L22 L30 0.298367
K22_31 L22 L31 0.015005
K22_32 L22 L32 0.0197607
K22_33 L22 L33 0.02423
K22_34 L22 L34 0.0276168
K22_35 L22 L35 0.0358181
K22_36 L22 L36 0.0198115
K22_37 L22 L37 -0.000237695
K22_38 L22 L38 -0.0183105
K23_24 L23 L24 0.941676
K23_25 L23 L25 0.879306
K23_26 L23 L26 0.298563
K23_27 L23 L27 0.306928
K23_28 L23 L28 0.324198
K23_29 L23 L29 0.321224
K23_30 L23 L30 0.313781
K23_31 L23 L31 0.0169833
K23_32 L23 L32 0.0200341
K23_33 L23 L33 0.0223757
K23_34 L23 L34 0.0236561
K23_35 L23 L35 0.0246966
K23_36 L23 L36 0.0221631
K23_37 L23 L37 0.0055108
K23_38 L23 L38 -0.0127072
K24_25 L24 L25 0.933804
K24_26 L24 L26 0.289002
K24_27 L24 L27 0.297145
K24_28 L24 L28 0.313881
K24_29 L24 L29 0.33346
K24_30 L24 L30 0.331497
K24_31 L24 L31 0.0196066
K24_32 L24 L32 0.0199425
K24_33 L24 L33 0.0197969
K24_34 L24 L34 0.0193924
K24_35 L24 L35 0.0147342
K24_36 L24 L36 0.0143891
K24_37 L24 L37 0.0122137
K24_38 L24 L38 -0.0021915
K25_26 L25 L26 0.276716
K25_27 L25 L27 0.284729
K25_28 L25 L28 0.30085
K25_29 L25 L29 0.319658
K25_30 L25 L30 0.343622
K25_31 L25 L31 0.0221394
K25_32 L25 L32 0.0197333
K25_33 L25 L33 0.017766
K25_34 L25 L34 0.0162614
K25_35 L25 L35 0.00814622
K25_36 L25 L36 0.00831304
K25_37 L25 L37 0.00879789
K25_38 L25 L38 0.0104079
K26_27 L26 L27 0.976612
K26_28 L26 L28 0.925223
K26_29 L26 L29 0.870316
K26_30 L26 L30 0.812315
K26_31 L26 L31 0.0120449
K26_32 L26 L32 0.0184609
K26_33 L26 L33 0.0244744
K26_34 L26 L34 0.0296343
K26_35 L26 L35 0.0272178
K26_36 L26 L36 0.0111498
K26_37 L26 L37 -0.00593148
K26_38 L26 L38 -0.0221974
K27_28 L27 L28 0.947533
K27_29 L27 L29 0.891284
K27_30 L27 L30 0.832066
K27_31 L27 L31 0.0144039
K27_32 L27 L32 0.0202608
K27_33 L27 L33 0.0255183
K27_34 L27 L34 0.0297238
K27_35 L27 L35 0.0289131
K27_36 L27 L36 0.014611
K27_37 L27 L37 -0.00238344
K27_38 L27 L38 -0.0188275
K28_29 L28 L29 0.941296
K28_30 L28 L30 0.878723
K28_31 L28 L31 0.0160516
K28_32 L28 L32 0.020601
K28_33 L28 L33 0.0241856
K28_34 L28 L34 0.0266099
K28_35 L28 L35 0.0227725
K28_36 L28 L36 0.0170063
K28_37 L28 L37 0.00181923
K28_38 L28 L38 -0.0147647
K29_30 L29 L30 0.933986
K29_31 L29 L31 0.0184534
K29_32 L29 L32 0.020817
K29_33 L29 L33 0.0222438
K29_34 L29 L34 0.023021
K29_35 L29 L35 0.0163037
K29_36 L29 L36 0.0145638
K29_37 L29 L37 0.00839928
K29_38 L29 L38 -0.00624289
K30_31 L30 L31 0.0210733
K30_32 L30 L32 0.0210069
K30_33 L30 L33 0.0206212
K30_34 L30 L34 0.0202226
K30_35 L30 L35 0.0123988
K30_36 L30 L36 0.0116076
K30_37 L30 L37 0.00989485
K30_38 L30 L38 0.00512309
K31_32 L31 L32 0.788974
K31_33 L31 L33 0.743965
K31_34 L31 L34 0.707954
K31_35 L31 L35 0.720366
K31_36 L31 L36 0.734832
K31_37 L31 L37 0.746384
K31_38 L31 L38 0.751767
K32_33 L32 L33 0.808835
K32_34 L32 L34 0.767478
K32_35 L32 L35 0.704641
K32_36 L32 L36 0.716271
K32_37 L32 L37 0.723083
K32_38 L32 L38 0.723784
K33_34 L33 L34 0.826439
K33_35 L33 L35 0.688166
K33_36 L33 L36 0.695651
K33_37 L33 L37 0.697887
K33_38 L33 L38 0.696002
K34_35 L34 L35 0.6696
K34_36 L34 L36 0.672567
K34_37 L34 L37 0.672022
K34_38 L34 L38 0.66881
K35_36 L35 L36 0.975796
K35_37 L35 L37 0.951012
K35_38 L35 L38 0.92539
K36_37 L36 L37 0.975051
K36_38 L36 L38 0.949233
K37_38 L37 L38 0.974278
.ends Quadraat_0004__4_0_4_0_4_0_4_half

.subckt Quadraat_0004__4_0_4_0_4_0_4_parlel 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15
+ 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38
C1_0 1 0 6.20836254827e-12
C1_5 1 5 3.23774759518e-15
C1_6 1 6 3.23774759518e-15
C1_7 1 7 3.23774759518e-15
C1_8 1 8 3.23774759518e-15
C1_9 1 9 3.23774759518e-15
C1_10 1 10 3.23774759518e-15
C1_11 1 11 3.23774759518e-15
C1_12 1 12 3.23774759518e-15
C1_13 1 13 3.23774759518e-15
C1_14 1 14 3.23774759518e-15
C1_15 1 15 3.23774759518e-15
C1_16 1 16 3.23774759518e-15
C1_17 1 17 3.23774759518e-15
C1_18 1 18 2.72700376666e-16
C1_19 1 19 2.03322622847e-16
C1_20 1 20 1.47690471994e-16
C1_21 1 21 1.08638587921e-16
C1_22 1 22 3.46007085613e-16
C1_23 1 23 3.46007085613e-16
C1_24 1 24 3.46007085613e-16
C1_25 1 25 3.46007085613e-16
C1_26 1 26 3.86552431369e-16
C1_27 1 27 3.86552431369e-16
C1_28 1 28 3.86552431369e-16
C1_29 1 29 3.86552431369e-16
C1_30 1 30 3.86552431369e-16
C1_31 1 31 6.06906228818e-13
C1_32 1 32 6.06906228818e-13
C1_33 1 33 6.06906228818e-13
C1_34 1 34 6.06906228818e-13
C1_35 1 35 6.06906228818e-13
C1_36 1 36 6.06906228818e-13
C1_37 1 37 6.06906228818e-13
C1_38 1 38 6.06906228818e-13
C2_0 2 0 6.20836254827e-12
C2_5 2 5 3.23774759518e-15
C2_6 2 6 3.23774759518e-15
C2_7 2 7 3.23774759518e-15
C2_8 2 8 3.23774759518e-15
C2_9 2 9 3.23774759518e-15
C2_10 2 10 3.23774759518e-15
C2_11 2 11 3.23774759518e-15
C2_12 2 12 3.23774759518e-15
C2_13 2 13 3.23774759518e-15
C2_14 2 14 3.23774759518e-15
C2_15 2 15 3.23774759518e-15
C2_16 2 16 3.23774759518e-15
C2_17 2 17 3.23774759518e-15
C2_18 2 18 2.72700376666e-16
C2_19 2 19 2.03322622847e-16
C2_20 2 20 1.47690471994e-16
C2_21 2 21 1.08638587921e-16
C2_22 2 22 3.46007085613e-16
C2_23 2 23 3.46007085613e-16
C2_24 2 24 3.46007085613e-16
C2_25 2 25 3.46007085613e-16
C2_26 2 26 3.86552431369e-16
C2_27 2 27 3.86552431369e-16
C2_28 2 28 3.86552431369e-16
C2_29 2 29 3.86552431369e-16
C2_30 2 30 3.86552431369e-16
C2_31 2 31 6.06906228818e-13
C2_32 2 32 6.06906228818e-13
C2_33 2 33 6.06906228818e-13
C2_34 2 34 6.06906228818e-13
C2_35 2 35 6.06906228818e-13
C2_36 2 36 6.06906228818e-13
C2_37 2 37 6.06906228818e-13
C2_38 2 38 6.06906228818e-13
C3_0 3 0 6.20836254827e-12
C3_5 3 5 3.23774759518e-15
C3_6 3 6 3.23774759518e-15
C3_7 3 7 3.23774759518e-15
C3_8 3 8 3.23774759518e-15
C3_9 3 9 3.23774759518e-15
C3_10 3 10 3.23774759518e-15
C3_11 3 11 3.23774759518e-15
C3_12 3 12 3.23774759518e-15
C3_13 3 13 3.23774759518e-15
C3_14 3 14 3.23774759518e-15
C3_15 3 15 3.23774759518e-15
C3_16 3 16 3.23774759518e-15
C3_17 3 17 3.23774759518e-15
C3_18 3 18 2.72700376666e-16
C3_19 3 19 2.03322622847e-16
C3_20 3 20 1.47690471994e-16
C3_21 3 21 1.08638587921e-16
C3_22 3 22 3.46007085613e-16
C3_23 3 23 3.46007085613e-16
C3_24 3 24 3.46007085613e-16
C3_25 3 25 3.46007085613e-16
C3_26 3 26 3.86552431369e-16
C3_27 3 27 3.86552431369e-16
C3_28 3 28 3.86552431369e-16
C3_29 3 29 3.86552431369e-16
C3_30 3 30 3.86552431369e-16
C3_31 3 31 6.06906228818e-13
C3_32 3 32 6.06906228818e-13
C3_33 3 33 6.06906228818e-13
C3_34 3 34 6.06906228818e-13
C3_35 3 35 6.06906228818e-13
C3_36 3 36 6.06906228818e-13
C3_37 3 37 6.06906228818e-13
C3_38 3 38 6.06906228818e-13
C4_0 4 0 6.20836254827e-12
C4_5 4 5 3.23774759518e-15
C4_6 4 6 3.23774759518e-15
C4_7 4 7 3.23774759518e-15
C4_8 4 8 3.23774759518e-15
C4_9 4 9 3.23774759518e-15
C4_10 4 10 3.23774759518e-15
C4_11 4 11 3.23774759518e-15
C4_12 4 12 3.23774759518e-15
C4_13 4 13 3.23774759518e-15
C4_14 4 14 3.23774759518e-15
C4_15 4 15 3.23774759518e-15
C4_16 4 16 3.23774759518e-15
C4_17 4 17 3.23774759518e-15
C4_18 4 18 2.72700376666e-16
C4_19 4 19 2.03322622847e-16
C4_20 4 20 1.47690471994e-16
C4_21 4 21 1.08638587921e-16
C4_22 4 22 3.46007085613e-16
C4_23 4 23 3.46007085613e-16
C4_24 4 24 3.46007085613e-16
C4_25 4 25 3.46007085613e-16
C4_26 4 26 3.86552431369e-16
C4_27 4 27 3.86552431369e-16
C4_28 4 28 3.86552431369e-16
C4_29 4 29 3.86552431369e-16
C4_30 4 30 3.86552431369e-16
C4_31 4 31 6.06906228818e-13
C4_32 4 32 6.06906228818e-13
C4_33 4 33 6.06906228818e-13
C4_34 4 34 6.06906228818e-13
C4_35 4 35 6.06906228818e-13
C4_36 4 36 6.06906228818e-13
C4_37 4 37 6.06906228818e-13
C4_38 4 38 6.06906228818e-13
C5_0 5 0 2.27976464006e-12
C5_18 5 18 1.11673852316e-14
C5_19 5 19 1.09042312442e-14
C5_20 5 20 1.07914503195e-14
C5_21 5 21 1.03702198583e-14
C5_22 5 22 2.03806759705e-15
C5_23 5 23 2.03806759705e-15
C5_24 5 24 2.03806759705e-15
C5_25 5 25 2.03806759705e-15
C5_26 5 26 1.18080588856e-13
C5_27 5 27 1.18080588856e-13
C5_28 5 28 1.18080588856e-13
C5_29 5 29 1.18080588856e-13
C5_30 5 30 1.18080588856e-13
C5_31 5 31 1.086330221e-13
C5_32 5 32 1.086330221e-13
C5_33 5 33 1.086330221e-13
C5_34 5 34 1.086330221e-13
C5_35 5 35 1.086330221e-13
C5_36 5 36 1.086330221e-13
C5_37 5 37 1.086330221e-13
C5_38 5 38 1.086330221e-13
C6_0 6 0 2.27976464006e-12
C6_18 6 18 1.11673852316e-14
C6_19 6 19 1.09042312442e-14
C6_20 6 20 1.07914503195e-14
C6_21 6 21 1.03702198583e-14
C6_22 6 22 2.03806759705e-15
C6_23 6 23 2.03806759705e-15
C6_24 6 24 2.03806759705e-15
C6_25 6 25 2.03806759705e-15
C6_26 6 26 1.18080588856e-13
C6_27 6 27 1.18080588856e-13
C6_28 6 28 1.18080588856e-13
C6_29 6 29 1.18080588856e-13
C6_30 6 30 1.18080588856e-13
C6_31 6 31 1.086330221e-13
C6_32 6 32 1.086330221e-13
C6_33 6 33 1.086330221e-13
C6_34 6 34 1.086330221e-13
C6_35 6 35 1.086330221e-13
C6_36 6 36 1.086330221e-13
C6_37 6 37 1.086330221e-13
C6_38 6 38 1.086330221e-13
C7_0 7 0 2.27976464006e-12
C7_18 7 18 1.11673852316e-14
C7_19 7 19 1.09042312442e-14
C7_20 7 20 1.07914503195e-14
C7_21 7 21 1.03702198583e-14
C7_22 7 22 2.03806759705e-15
C7_23 7 23 2.03806759705e-15
C7_24 7 24 2.03806759705e-15
C7_25 7 25 2.03806759705e-15
C7_26 7 26 1.18080588856e-13
C7_27 7 27 1.18080588856e-13
C7_28 7 28 1.18080588856e-13
C7_29 7 29 1.18080588856e-13
C7_30 7 30 1.18080588856e-13
C7_31 7 31 1.086330221e-13
C7_32 7 32 1.086330221e-13
C7_33 7 33 1.086330221e-13
C7_34 7 34 1.086330221e-13
C7_35 7 35 1.086330221e-13
C7_36 7 36 1.086330221e-13
C7_37 7 37 1.086330221e-13
C7_38 7 38 1.086330221e-13
C8_0 8 0 2.27976464006e-12
C8_18 8 18 1.11673852316e-14
C8_19 8 19 1.09042312442e-14
C8_20 8 20 1.07914503195e-14
C8_21 8 21 1.03702198583e-14
C8_22 8 22 2.03806759705e-15
C8_23 8 23 2.03806759705e-15
C8_24 8 24 2.03806759705e-15
C8_25 8 25 2.03806759705e-15
C8_26 8 26 1.18080588856e-13
C8_27 8 27 1.18080588856e-13
C8_28 8 28 1.18080588856e-13
C8_29 8 29 1.18080588856e-13
C8_30 8 30 1.18080588856e-13
C8_31 8 31 1.086330221e-13
C8_32 8 32 1.086330221e-13
C8_33 8 33 1.086330221e-13
C8_34 8 34 1.086330221e-13
C8_35 8 35 1.086330221e-13
C8_36 8 36 1.086330221e-13
C8_37 8 37 1.086330221e-13
C8_38 8 38 1.086330221e-13
C9_0 9 0 2.27976464006e-12
C9_18 9 18 1.11673852316e-14
C9_19 9 19 1.09042312442e-14
C9_20 9 20 1.07914503195e-14
C9_21 9 21 1.03702198583e-14
C9_22 9 22 2.03806759705e-15
C9_23 9 23 2.03806759705e-15
C9_24 9 24 2.03806759705e-15
C9_25 9 25 2.03806759705e-15
C9_26 9 26 1.18080588856e-13
C9_27 9 27 1.18080588856e-13
C9_28 9 28 1.18080588856e-13
C9_29 9 29 1.18080588856e-13
C9_30 9 30 1.18080588856e-13
C9_31 9 31 1.086330221e-13
C9_32 9 32 1.086330221e-13
C9_33 9 33 1.086330221e-13
C9_34 9 34 1.086330221e-13
C9_35 9 35 1.086330221e-13
C9_36 9 36 1.086330221e-13
C9_37 9 37 1.086330221e-13
C9_38 9 38 1.086330221e-13
C10_0 10 0 2.27976464006e-12
C10_18 10 18 1.11673852316e-14
C10_19 10 19 1.09042312442e-14
C10_20 10 20 1.07914503195e-14
C10_21 10 21 1.03702198583e-14
C10_22 10 22 2.03806759705e-15
C10_23 10 23 2.03806759705e-15
C10_24 10 24 2.03806759705e-15
C10_25 10 25 2.03806759705e-15
C10_26 10 26 1.18080588856e-13
C10_27 10 27 1.18080588856e-13
C10_28 10 28 1.18080588856e-13
C10_29 10 29 1.18080588856e-13
C10_30 10 30 1.18080588856e-13
C10_31 10 31 1.086330221e-13
C10_32 10 32 1.086330221e-13
C10_33 10 33 1.086330221e-13
C10_34 10 34 1.086330221e-13
C10_35 10 35 1.086330221e-13
C10_36 10 36 1.086330221e-13
C10_37 10 37 1.086330221e-13
C10_38 10 38 1.086330221e-13
C11_0 11 0 2.27976464006e-12
C11_18 11 18 1.11673852316e-14
C11_19 11 19 1.09042312442e-14
C11_20 11 20 1.07914503195e-14
C11_21 11 21 1.03702198583e-14
C11_22 11 22 2.03806759705e-15
C11_23 11 23 2.03806759705e-15
C11_24 11 24 2.03806759705e-15
C11_25 11 25 2.03806759705e-15
C11_26 11 26 1.18080588856e-13
C11_27 11 27 1.18080588856e-13
C11_28 11 28 1.18080588856e-13
C11_29 11 29 1.18080588856e-13
C11_30 11 30 1.18080588856e-13
C11_31 11 31 1.086330221e-13
C11_32 11 32 1.086330221e-13
C11_33 11 33 1.086330221e-13
C11_34 11 34 1.086330221e-13
C11_35 11 35 1.086330221e-13
C11_36 11 36 1.086330221e-13
C11_37 11 37 1.086330221e-13
C11_38 11 38 1.086330221e-13
C12_0 12 0 2.27976464006e-12
C12_18 12 18 1.11673852316e-14
C12_19 12 19 1.09042312442e-14
C12_20 12 20 1.07914503195e-14
C12_21 12 21 1.03702198583e-14
C12_22 12 22 2.03806759705e-15
C12_23 12 23 2.03806759705e-15
C12_24 12 24 2.03806759705e-15
C12_25 12 25 2.03806759705e-15
C12_26 12 26 1.18080588856e-13
C12_27 12 27 1.18080588856e-13
C12_28 12 28 1.18080588856e-13
C12_29 12 29 1.18080588856e-13
C12_30 12 30 1.18080588856e-13
C12_31 12 31 1.086330221e-13
C12_32 12 32 1.086330221e-13
C12_33 12 33 1.086330221e-13
C12_34 12 34 1.086330221e-13
C12_35 12 35 1.086330221e-13
C12_36 12 36 1.086330221e-13
C12_37 12 37 1.086330221e-13
C12_38 12 38 1.086330221e-13
C13_0 13 0 2.27976464006e-12
C13_18 13 18 1.11673852316e-14
C13_19 13 19 1.09042312442e-14
C13_20 13 20 1.07914503195e-14
C13_21 13 21 1.03702198583e-14
C13_22 13 22 2.03806759705e-15
C13_23 13 23 2.03806759705e-15
C13_24 13 24 2.03806759705e-15
C13_25 13 25 2.03806759705e-15
C13_26 13 26 1.18080588856e-13
C13_27 13 27 1.18080588856e-13
C13_28 13 28 1.18080588856e-13
C13_29 13 29 1.18080588856e-13
C13_30 13 30 1.18080588856e-13
C13_31 13 31 1.086330221e-13
C13_32 13 32 1.086330221e-13
C13_33 13 33 1.086330221e-13
C13_34 13 34 1.086330221e-13
C13_35 13 35 1.086330221e-13
C13_36 13 36 1.086330221e-13
C13_37 13 37 1.086330221e-13
C13_38 13 38 1.086330221e-13
C14_0 14 0 2.27976464006e-12
C14_18 14 18 1.11673852316e-14
C14_19 14 19 1.09042312442e-14
C14_20 14 20 1.07914503195e-14
C14_21 14 21 1.03702198583e-14
C14_22 14 22 2.03806759705e-15
C14_23 14 23 2.03806759705e-15
C14_24 14 24 2.03806759705e-15
C14_25 14 25 2.03806759705e-15
C14_26 14 26 1.18080588856e-13
C14_27 14 27 1.18080588856e-13
C14_28 14 28 1.18080588856e-13
C14_29 14 29 1.18080588856e-13
C14_30 14 30 1.18080588856e-13
C14_31 14 31 1.086330221e-13
C14_32 14 32 1.086330221e-13
C14_33 14 33 1.086330221e-13
C14_34 14 34 1.086330221e-13
C14_35 14 35 1.086330221e-13
C14_36 14 36 1.086330221e-13
C14_37 14 37 1.086330221e-13
C14_38 14 38 1.086330221e-13
C15_0 15 0 2.27976464006e-12
C15_18 15 18 1.11673852316e-14
C15_19 15 19 1.09042312442e-14
C15_20 15 20 1.07914503195e-14
C15_21 15 21 1.03702198583e-14
C15_22 15 22 2.03806759705e-15
C15_23 15 23 2.03806759705e-15
C15_24 15 24 2.03806759705e-15
C15_25 15 25 2.03806759705e-15
C15_26 15 26 1.18080588856e-13
C15_27 15 27 1.18080588856e-13
C15_28 15 28 1.18080588856e-13
C15_29 15 29 1.18080588856e-13
C15_30 15 30 1.18080588856e-13
C15_31 15 31 1.086330221e-13
C15_32 15 32 1.086330221e-13
C15_33 15 33 1.086330221e-13
C15_34 15 34 1.086330221e-13
C15_35 15 35 1.086330221e-13
C15_36 15 36 1.086330221e-13
C15_37 15 37 1.086330221e-13
C15_38 15 38 1.086330221e-13
C16_0 16 0 2.27976464006e-12
C16_18 16 18 1.11673852316e-14
C16_19 16 19 1.09042312442e-14
C16_20 16 20 1.07914503195e-14
C16_21 16 21 1.03702198583e-14
C16_22 16 22 2.03806759705e-15
C16_23 16 23 2.03806759705e-15
C16_24 16 24 2.03806759705e-15
C16_25 16 25 2.03806759705e-15
C16_26 16 26 1.18080588856e-13
C16_27 16 27 1.18080588856e-13
C16_28 16 28 1.18080588856e-13
C16_29 16 29 1.18080588856e-13
C16_30 16 30 1.18080588856e-13
C16_31 16 31 1.086330221e-13
C16_32 16 32 1.086330221e-13
C16_33 16 33 1.086330221e-13
C16_34 16 34 1.086330221e-13
C16_35 16 35 1.086330221e-13
C16_36 16 36 1.086330221e-13
C16_37 16 37 1.086330221e-13
C16_38 16 38 1.086330221e-13
C17_0 17 0 2.27976464006e-12
C17_18 17 18 1.11673852316e-14
C17_19 17 19 1.09042312442e-14
C17_20 17 20 1.07914503195e-14
C17_21 17 21 1.03702198583e-14
C17_22 17 22 2.03806759705e-15
C17_23 17 23 2.03806759705e-15
C17_24 17 24 2.03806759705e-15
C17_25 17 25 2.03806759705e-15
C17_26 17 26 1.18080588856e-13
C17_27 17 27 1.18080588856e-13
C17_28 17 28 1.18080588856e-13
C17_29 17 29 1.18080588856e-13
C17_30 17 30 1.18080588856e-13
C17_31 17 31 1.086330221e-13
C17_32 17 32 1.086330221e-13
C17_33 17 33 1.086330221e-13
C17_34 17 34 1.086330221e-13
C17_35 17 35 1.086330221e-13
C17_36 17 36 1.086330221e-13
C17_37 17 37 1.086330221e-13
C17_38 17 38 1.086330221e-13
C18_0 18 0 2.92365892259e-14
C18_19 18 19 1.05814590562e-15
C18_20 18 20 1.60915761221e-16
C18_21 18 21 4.81605481136e-17
C18_22 18 22 4.71320970215e-13
C18_23 18 23 4.71320970215e-13
C18_24 18 24 4.71320970215e-13
C18_25 18 25 4.71320970215e-13
C18_26 18 26 3.12860445446e-15
C18_27 18 27 3.12860445446e-15
C18_28 18 28 3.12860445446e-15
C18_29 18 29 3.12860445446e-15
C18_30 18 30 3.12860445446e-15
C18_31 18 31 7.11700978363e-14
C18_32 18 32 7.11700978363e-14
C18_33 18 33 7.11700978363e-14
C18_34 18 34 7.11700978363e-14
C18_35 18 35 7.11700978363e-14
C18_36 18 36 7.11700978363e-14
C18_37 18 37 7.11700978363e-14
C18_38 18 38 7.11700978363e-14
C19_0 19 0 2.9393335868e-14
C19_20 19 20 1.07304460083e-15
C19_21 19 21 1.36760340994e-16
C19_22 19 22 4.72130735851e-13
C19_23 19 23 4.72130735851e-13
C19_24 19 24 4.72130735851e-13
C19_25 19 25 4.72130735851e-13
C19_26 19 26 2.71522992467e-15
C19_27 19 27 2.71522992467e-15
C19_28 19 28 2.71522992467e-15
C19_29 19 29 2.71522992467e-15
C19_30 19 30 2.71522992467e-15
C19_31 19 31 7.12960754523e-14
C19_32 19 32 7.12960754523e-14
C19_33 19 33 7.12960754523e-14
C19_34 19 34 7.12960754523e-14
C19_35 19 35 7.12960754523e-14
C19_36 19 36 7.12960754523e-14
C19_37 19 37 7.12960754523e-14
C19_38 19 38 7.12960754523e-14
C20_0 20 0 2.83967273964e-14
C20_21 20 21 9.81388407004e-16
C20_22 20 22 4.72577207422e-13
C20_23 20 23 4.72577207422e-13
C20_24 20 24 4.72577207422e-13
C20_25 20 25 4.72577207422e-13
C20_26 20 26 2.7351613348e-15
C20_27 20 27 2.7351613348e-15
C20_28 20 28 2.7351613348e-15
C20_29 20 29 2.7351613348e-15
C20_30 20 30 2.7351613348e-15
C20_31 20 31 7.13213387428e-14
C20_32 20 32 7.13213387428e-14
C20_33 20 33 7.13213387428e-14
C20_34 20 34 7.13213387428e-14
C20_35 20 35 7.13213387428e-14
C20_36 20 36 7.13213387428e-14
C20_37 20 37 7.13213387428e-14
C20_38 20 38 7.13213387428e-14
C21_0 21 0 2.86880202781e-14
C21_22 21 22 4.74599604762e-13
C21_23 21 23 4.74599604762e-13
C21_24 21 24 4.74599604762e-13
C21_25 21 25 4.74599604762e-13
C21_26 21 26 2.85622166275e-15
C21_27 21 27 2.85622166275e-15
C21_28 21 28 2.85622166275e-15
C21_29 21 29 2.85622166275e-15
C21_30 21 30 2.85622166275e-15
C21_31 21 31 7.11415025923e-14
C21_32 21 32 7.11415025923e-14
C21_33 21 33 7.11415025923e-14
C21_34 21 34 7.11415025923e-14
C21_35 21 35 7.11415025923e-14
C21_36 21 36 7.11415025923e-14
C21_37 21 37 7.11415025923e-14
C21_38 21 38 7.11415025923e-14
C22_0 22 0 1.60239003518e-12
C22_26 22 26 6.98489999477e-14
C22_27 22 27 6.98489999477e-14
C22_28 22 28 6.98489999477e-14
C22_29 22 29 6.98489999477e-14
C22_30 22 30 6.98489999477e-14
C22_31 22 31 1.06789200723e-14
C22_32 22 32 1.06789200723e-14
C22_33 22 33 1.06789200723e-14
C22_34 22 34 1.06789200723e-14
C22_35 22 35 1.06789200723e-14
C22_36 22 36 1.06789200723e-14
C22_37 22 37 1.06789200723e-14
C22_38 22 38 1.06789200723e-14
C23_0 23 0 1.60239003518e-12
C23_26 23 26 6.98489999477e-14
C23_27 23 27 6.98489999477e-14
C23_28 23 28 6.98489999477e-14
C23_29 23 29 6.98489999477e-14
C23_30 23 30 6.98489999477e-14
C23_31 23 31 1.06789200723e-14
C23_32 23 32 1.06789200723e-14
C23_33 23 33 1.06789200723e-14
C23_34 23 34 1.06789200723e-14
C23_35 23 35 1.06789200723e-14
C23_36 23 36 1.06789200723e-14
C23_37 23 37 1.06789200723e-14
C23_38 23 38 1.06789200723e-14
C24_0 24 0 1.60239003518e-12
C24_26 24 26 6.98489999477e-14
C24_27 24 27 6.98489999477e-14
C24_28 24 28 6.98489999477e-14
C24_29 24 29 6.98489999477e-14
C24_30 24 30 6.98489999477e-14
C24_31 24 31 1.06789200723e-14
C24_32 24 32 1.06789200723e-14
C24_33 24 33 1.06789200723e-14
C24_34 24 34 1.06789200723e-14
C24_35 24 35 1.06789200723e-14
C24_36 24 36 1.06789200723e-14
C24_37 24 37 1.06789200723e-14
C24_38 24 38 1.06789200723e-14
C25_0 25 0 1.60239003518e-12
C25_26 25 26 6.98489999477e-14
C25_27 25 27 6.98489999477e-14
C25_28 25 28 6.98489999477e-14
C25_29 25 29 6.98489999477e-14
C25_30 25 30 6.98489999477e-14
C25_31 25 31 1.06789200723e-14
C25_32 25 32 1.06789200723e-14
C25_33 25 33 1.06789200723e-14
C25_34 25 34 1.06789200723e-14
C25_35 25 35 1.06789200723e-14
C25_36 25 36 1.06789200723e-14
C25_37 25 37 1.06789200723e-14
C25_38 25 38 1.06789200723e-14
C26_0 26 0 1.48209127357e-12
C26_31 26 31 2.14588123681e-15
C26_32 26 32 2.14588123681e-15
C26_33 26 33 2.14588123681e-15
C26_34 26 34 2.14588123681e-15
C26_35 26 35 2.14588123681e-15
C26_36 26 36 2.14588123681e-15
C26_37 26 37 2.14588123681e-15
C26_38 26 38 2.14588123681e-15
C27_0 27 0 1.48209127357e-12
C27_31 27 31 2.14588123681e-15
C27_32 27 32 2.14588123681e-15
C27_33 27 33 2.14588123681e-15
C27_34 27 34 2.14588123681e-15
C27_35 27 35 2.14588123681e-15
C27_36 27 36 2.14588123681e-15
C27_37 27 37 2.14588123681e-15
C27_38 27 38 2.14588123681e-15
C28_0 28 0 1.48209127357e-12
C28_31 28 31 2.14588123681e-15
C28_32 28 32 2.14588123681e-15
C28_33 28 33 2.14588123681e-15
C28_34 28 34 2.14588123681e-15
C28_35 28 35 2.14588123681e-15
C28_36 28 36 2.14588123681e-15
C28_37 28 37 2.14588123681e-15
C28_38 28 38 2.14588123681e-15
C29_0 29 0 1.48209127357e-12
C29_31 29 31 2.14588123681e-15
C29_32 29 32 2.14588123681e-15
C29_33 29 33 2.14588123681e-15
C29_34 29 34 2.14588123681e-15
C29_35 29 35 2.14588123681e-15
C29_36 29 36 2.14588123681e-15
C29_37 29 37 2.14588123681e-15
C29_38 29 38 2.14588123681e-15
C30_0 30 0 1.48209127357e-12
C30_31 30 31 2.14588123681e-15
C30_32 30 32 2.14588123681e-15
C30_33 30 33 2.14588123681e-15
C30_34 30 34 2.14588123681e-15
C30_35 30 35 2.14588123681e-15
C30_36 30 36 2.14588123681e-15
C30_37 30 37 2.14588123681e-15
C30_38 30 38 2.14588123681e-15
C31_0 31 0 7.59590584832e-12
C32_0 32 0 7.59590584832e-12
C33_0 33 0 7.59590584832e-12
C34_0 34 0 7.59590584832e-12
C35_0 35 0 7.59590584832e-12
C36_0 36 0 7.59590584832e-12
C37_0 37 0 7.59590584832e-12
C38_0 38 0 7.59590584832e-12
.ends Quadraat_0004__4_0_4_0_4_0_4_parlel

.ends Quadraat_0004__4_0_4_0_4_0_4
