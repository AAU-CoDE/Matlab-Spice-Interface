* BEGIN ANSOFT HEADER
* node 1    DC+:D1K
* node 2    DC+:D2K
* node 3    DC+:D3K
* node 4    DC+:D4K
* node 5    DC-:DC-GS-short-b
* node 6    DC-:Q1BW
* node 7    DC-:Q1S
* node 8    DC-:Q2BW
* node 9    DC-:Q2S
* node 10   DC-:Q3BW
* node 11   DC-:Q3S
* node 12   DC-:Q4BW
* node 13   DC-:Q4S
* node 14   DC-:RS1b
* node 15   DC-:RS2b
* node 16   DC-:RS3b
* node 17   DC-:RS4b
* node 18   G1:Q1G
* node 19   G2:Q2G
* node 20   G3:Q3G
* node 21   G4:Q4G
* node 22   GG:RG1a
* node 23   GG:RG2a
* node 24   GG:RG3a
* node 25   GG:RG4a
* node 26   GS:DC-GS-short-a
* node 27   GS:RS1a
* node 28   GS:RS2a
* node 29   GS:RS3a
* node 30   GS:RS4a
* node 31   OUT:D1A
* node 32   OUT:D2A
* node 33   OUT:D3A
* node 34   OUT:D4A
* node 35   OUT:Q1D
* node 36   OUT:Q2D
* node 37   OUT:Q3D
* node 38   OUT:Q4D
* node 39   DC+:DC+terminal
* node 40   DC-:DC-terminal
* node 41   G1:RG1b
* node 42   G2:RG2b
* node 43   G3:RG3b
* node 44   G4:RG4b
* node 45   GG:G-terminal
* node 46   GS:S-terminal
* node 47   OUT:OUT-terminal
*  Project: Quadraat 0004 [7.0 6.0 5.0 4.0]
*   Design: Q3DDesign1
*   Format: Ansys Nexxim
*   Topckt: Quadraat_0004__7_0_6_0_5_0_4
*  Creator: Ansys Electronics Desktop 2022.1.0
*     Date: Wed Nov 30 15:12:00 2022
* END ANSOFT HEADER

.subckt Quadraat 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17
+ 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42 43
+ 44 45 46 47
X1 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29
+ 30 31 32 33 34 35 36 37 38 39 39 39 39 40 40 40 40 40 40 40 40 40 40 40 40 40
+ 41 42 43 44 45 45 45 45 46 46 46 46 46 47 47 47 47 47 47 47 47
+ Quadraat_0004__7_0_6_0_5_0_4_series

.subckt Quadraat_0004__7_0_6_0_5_0_4_series 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15
+ 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41
+ 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62 63 64 65 66 67
+ 68 69 70 71 72 73 74 75 76
V1 1 77 dc 0.0
V2 2 78 dc 0.0
V3 3 79 dc 0.0
V4 4 80 dc 0.0
V5 5 81 dc 0.0
V6 6 82 dc 0.0
V7 7 83 dc 0.0
V8 8 84 dc 0.0
V9 9 85 dc 0.0
V10 10 86 dc 0.0
V11 11 87 dc 0.0
V12 12 88 dc 0.0
V13 13 89 dc 0.0
V14 14 90 dc 0.0
V15 15 91 dc 0.0
V16 16 92 dc 0.0
V17 17 93 dc 0.0
V18 18 94 dc 0.0
V19 19 95 dc 0.0
V20 20 96 dc 0.0
V21 21 97 dc 0.0
V22 22 98 dc 0.0
V23 23 99 dc 0.0
V24 24 100 dc 0.0
V25 25 101 dc 0.0
V26 26 102 dc 0.0
V27 27 103 dc 0.0
V28 28 104 dc 0.0
V29 29 105 dc 0.0
V30 30 106 dc 0.0
V31 31 107 dc 0.0
V32 32 108 dc 0.0
V33 33 109 dc 0.0
V34 34 110 dc 0.0
V35 35 111 dc 0.0
V36 36 112 dc 0.0
V37 37 113 dc 0.0
V38 38 114 dc 0.0
R1 77 115 0.00102177046678
R2 78 116 0.000975131183416
R3 79 117 0.000928229437958
R4 80 118 0.00088170252132
R5 81 119 0.00159968719842
R6 82 120 0.000985279468314
R7 83 121 0.00322533520483
R8 84 122 0.00107052895838
R9 85 123 0.00306632737961
R10 86 124 0.00115196700505
R11 87 125 0.00293835515515
R12 88 126 0.00124267499614
R13 89 127 0.0028361533485
R14 90 128 0.00720314461879
R15 91 129 0.00704615368808
R16 92 130 0.00692684427475
R17 93 131 0.00680831719631
R18 94 132 0.00366611434531
R19 95 133 0.00365432708298
R20 96 134 0.00365491262192
R21 97 135 0.00366302058211
R22 98 136 0.00502915936896
R23 99 137 0.00462608842597
R24 100 138 0.00422197249329
R25 101 139 0.00381840211701
R26 102 140 0.00541729772822
R27 103 141 0.00465760625101
R28 104 142 0.00425550231535
R29 105 143 0.00385367932913
R30 106 144 0.00345325029543
R31 107 145 0.00314383156312
R32 108 146 0.003267333718
R33 109 147 0.00339138960373
R34 110 148 0.00350992867179
R35 111 149 0.00185284563642
R36 112 150 0.00180799080012
R37 113 151 0.00176343888287
R38 114 152 0.00171969500213
F1_2 115 77 V2 0.95401
F1_3 115 77 V3 0.90814
F1_4 115 77 V4 0.862632
F2_1 116 78 V1 0.999639
F2_3 116 78 V3 0.951575
F2_4 116 78 V4 0.903891
F3_1 117 79 V1 0.999656
F3_2 117 79 V2 0.999656
F3_4 117 79 V4 0.949563
F4_1 118 80 V1 0.999671
F4_2 118 80 V2 0.999671
F4_3 118 80 V3 0.999671
F5_6 119 81 V6 0.512946
F5_7 119 81 V7 0.512946
F5_8 119 81 V8 0.512946
F5_9 119 81 V9 0.512946
F5_10 119 81 V10 0.512946
F5_11 119 81 V11 0.512946
F5_12 119 81 V12 0.512946
F5_13 119 81 V13 0.512946
F5_14 119 81 V14 0.512946
F5_15 119 81 V15 0.512946
F5_16 119 81 V16 0.512946
F5_17 119 81 V17 0.512946
F6_5 120 82 V5 0.832812
F6_7 120 82 V7 0.992443
F6_8 120 82 V8 0.987844
F6_9 120 82 V9 0.987822
F6_10 120 82 V10 0.987842
F6_11 120 82 V11 0.987842
F6_12 120 82 V12 0.987842
F6_13 120 82 V13 0.987842
F6_14 120 82 V14 0.992443
F6_15 120 82 V15 0.987822
F6_16 120 82 V16 0.987842
F6_17 120 82 V17 0.987842
F7_5 121 83 V5 0.254409
F7_6 121 83 V6 0.303173
F7_8 121 83 V8 0.301805
F7_9 121 83 V9 0.3018
F7_10 121 83 V10 0.301804
F7_11 121 83 V11 0.301804
F7_12 121 83 V12 0.301804
F7_13 121 83 V13 0.301804
F7_14 121 83 V14 1.00003
F7_15 121 83 V15 0.3018
F7_16 121 83 V16 0.301804
F7_17 121 83 V17 0.301804
F8_5 122 84 V5 0.766494
F8_6 122 84 V6 0.909179
F8_7 122 84 V7 0.90929
F8_9 122 84 V9 0.989383
F8_10 122 84 V10 0.985269
F8_11 122 84 V11 0.985269
F8_12 122 84 V12 0.98527
F8_13 122 84 V13 0.98527
F8_14 122 84 V14 0.909291
F8_15 122 84 V15 0.989383
F8_16 122 84 V16 0.985269
F8_17 122 84 V17 0.98527
F9_5 123 85 V5 0.267601
F9_6 123 85 V6 0.317409
F9_7 123 85 V7 0.31745
F9_8 123 85 V8 0.345418
F9_10 123 85 V10 0.343942
F9_11 123 85 V11 0.343944
F9_12 123 85 V12 0.343936
F9_13 123 85 V13 0.343936
F9_14 123 85 V14 0.31745
F9_15 123 85 V15 1
F9_16 123 85 V16 0.343944
F9_17 123 85 V17 0.343936
F10_5 124 86 V5 0.712307
F10_6 124 86 V6 0.844903
F10_7 124 86 V7 0.845006
F10_8 124 86 V8 0.915616
F10_9 124 86 V9 0.915512
F10_11 124 86 V11 0.992647
F10_12 124 86 V12 0.986578
F10_13 124 86 V13 0.98658
F10_14 124 86 V14 0.845007
F10_15 124 86 V15 0.915512
F10_16 124 86 V16 0.992647
F10_17 124 86 V17 0.98658
F11_5 125 87 V5 0.279256
F11_6 125 87 V6 0.33124
F11_7 125 87 V7 0.33128
F11_8 125 87 V8 0.358962
F11_9 125 87 V9 0.358923
F11_10 125 87 V10 0.389162
F11_12 125 87 V12 0.386792
F11_13 125 87 V13 0.386792
F11_14 125 87 V14 0.33128
F11_15 125 87 V15 0.358923
F11_16 125 87 V16 1
F11_17 125 87 V17 0.386792
F12_5 126 88 V5 0.660312
F12_6 126 88 V6 0.78323
F12_7 126 88 V7 0.783326
F12_8 126 88 V8 0.848782
F12_9 126 88 V9 0.84867
F12_10 126 88 V10 0.914564
F12_11 126 88 V11 0.914584
F12_13 126 88 V13 0.997266
F12_14 126 88 V14 0.783326
F12_15 126 88 V15 0.84867
F12_16 126 88 V16 0.914584
F12_17 126 88 V17 0.997266
F13_5 127 89 V5 0.289319
F13_6 127 89 V6 0.343176
F13_7 127 89 V7 0.343218
F13_8 127 89 V8 0.371898
F13_9 127 89 V9 0.371849
F13_10 127 89 V10 0.400721
F13_11 127 89 V11 0.40073
F13_12 127 89 V12 0.436957
F13_14 127 89 V14 0.343218
F13_15 127 89 V15 0.371849
F13_16 127 89 V16 0.40073
F13_17 127 89 V17 1
F14_5 128 90 V5 0.113916
F14_6 128 90 V6 0.135751
F14_7 128 90 V7 0.447782
F14_8 128 90 V8 0.135138
F14_9 128 90 V9 0.135136
F14_10 128 90 V10 0.135138
F14_11 128 90 V11 0.135138
F14_12 128 90 V12 0.135138
F14_13 128 90 V13 0.135138
F14_15 128 90 V15 0.135136
F14_16 128 90 V16 0.135138
F14_17 128 90 V17 0.135138
F15_5 129 91 V5 0.116454
F15_6 129 91 V6 0.138129
F15_7 129 91 V7 0.138147
F15_8 129 91 V8 0.150318
F15_9 129 91 V9 0.435178
F15_10 129 91 V10 0.149676
F15_11 129 91 V11 0.149677
F15_12 129 91 V12 0.149673
F15_13 129 91 V13 0.149673
F15_14 129 91 V14 0.138147
F15_16 129 91 V16 0.149677
F15_17 129 91 V17 0.149673
F16_5 130 92 V5 0.11846
F16_6 130 92 V6 0.140511
F16_7 130 92 V7 0.140529
F16_8 130 92 V8 0.152271
F16_9 130 92 V9 0.152255
F16_10 130 92 V10 0.165082
F16_11 130 92 V11 0.424198
F16_12 130 92 V12 0.164076
F16_13 130 92 V13 0.164077
F16_14 130 92 V14 0.140529
F16_15 130 92 V15 0.152255
F16_17 130 92 V17 0.164077
F17_5 131 93 V5 0.120522
F17_6 131 93 V6 0.142958
F17_7 131 93 V7 0.142975
F17_8 131 93 V8 0.154922
F17_9 131 93 V9 0.154902
F17_10 131 93 V10 0.166929
F17_11 131 93 V11 0.166933
F17_12 131 93 V12 0.182024
F17_13 131 93 V13 0.416572
F17_14 131 93 V14 0.142975
F17_15 131 93 V15 0.154902
F17_16 131 93 V16 0.166933
F22_23 136 98 V23 0.919835
F22_24 136 98 V24 0.83948
F22_25 136 98 V25 0.759235
F23_22 137 99 V22 0.99998
F23_24 137 99 V24 0.912624
F23_25 137 99 V25 0.825387
F24_22 138 100 V22 0.999978
F24_23 138 100 V23 0.999978
F24_25 138 100 V25 0.904391
F25_22 139 101 V22 0.999977
F25_23 139 101 V23 0.999977
F25_24 139 101 V24 0.999977
F26_27 140 102 V27 0.85974
F26_28 140 102 V28 0.785524
F26_29 140 102 V29 0.711351
F26_30 140 102 V30 0.637436
F27_26 141 103 V26 0.99997
F27_28 141 103 V28 0.913649
F27_29 141 103 V29 0.827377
F27_30 141 103 V30 0.741407
F28_26 142 104 V26 0.99998
F28_27 142 104 V27 0.99998
F28_29 142 104 V29 0.905557
F28_30 142 104 V30 0.811463
F29_26 143 105 V26 0.999979
F29_27 143 105 V27 0.999979
F29_28 143 105 V28 0.999979
F29_30 143 105 V30 0.896074
F30_26 144 106 V26 0.99998
F30_27 144 106 V27 0.99998
F30_28 144 106 V28 0.99998
F30_29 144 106 V29 0.99998
F31_32 145 107 V32 0.492271
F31_33 145 107 V33 0.492256
F31_34 145 107 V34 0.492256
F31_35 145 107 V35 0.464483
F31_36 145 107 V36 0.464483
F31_37 145 107 V37 0.464483
F31_38 145 107 V38 0.464483
F32_31 146 108 V31 0.473664
F32_33 146 108 V33 0.511434
F32_34 146 108 V34 0.511435
F32_35 146 108 V35 0.446979
F32_36 146 108 V36 0.446979
F32_37 146 108 V37 0.446979
F32_38 146 108 V38 0.446979
F33_31 147 109 V31 0.456323
F33_32 147 109 V32 0.492726
F33_34 147 109 V34 0.528973
F33_35 147 109 V35 0.430631
F33_36 147 109 V36 0.430631
F33_37 147 109 V37 0.430631
F33_38 147 109 V38 0.430631
F34_31 148 110 V31 0.440912
F34_32 148 110 V32 0.476086
F34_33 148 110 V33 0.511108
F34_35 148 110 V35 0.416088
F34_36 148 110 V36 0.416088
F34_37 148 110 V37 0.416088
F34_38 148 110 V38 0.416088
F35_31 149 111 V31 0.788116
F35_32 149 111 V32 0.788209
F35_33 149 111 V33 0.788213
F35_34 149 111 V34 0.788213
F35_36 149 111 V36 0.975053
F35_37 149 111 V37 0.950997
F35_38 149 111 V38 0.927111
F36_31 150 112 V31 0.807669
F36_32 150 112 V32 0.807764
F36_33 150 112 V33 0.807768
F36_34 150 112 V34 0.807768
F36_35 150 112 V35 0.999243
F36_37 150 112 V37 0.974593
F36_38 150 112 V38 0.950112
F37_31 151 113 V31 0.828074
F37_32 151 113 V32 0.828172
F37_33 151 113 V33 0.828176
F37_34 151 113 V34 0.828176
F37_35 151 113 V35 0.999212
F37_36 151 113 V36 0.999215
F37_38 151 113 V38 0.974119
F38_31 152 114 V31 0.849137
F38_32 152 114 V32 0.849238
F38_33 152 114 V33 0.849242
F38_34 152 114 V34 0.849242
F38_35 152 114 V35 0.998895
F38_36 152 114 V36 0.998895
F38_37 152 114 V37 0.998898
L1 115 39 9.81357293772e-09
L2 116 40 9.14550153964e-09
L3 117 41 8.44830720146e-09
L4 118 42 7.67147115842e-09
L5 119 43 7.53735944938e-09
L6 120 44 9.2255737207e-09
L7 121 45 1.15177010479e-08
L8 122 46 1.02630310557e-08
L9 123 47 1.26704067083e-08
L10 124 48 1.13933937634e-08
L11 125 49 1.36835888346e-08
L12 126 50 1.26606025854e-08
L13 127 51 1.47519056472e-08
L14 128 52 1.53489728021e-08
L15 129 53 1.66155424013e-08
L16 130 54 1.76683005079e-08
L17 131 55 1.87587182958e-08
L18 132 56 3.63720655108e-09
L19 133 57 3.63244843786e-09
L20 134 58 3.63317703234e-09
L21 135 59 3.65236972998e-09
L22 136 60 1.56137961302e-08
L23 137 61 1.40090532241e-08
L24 138 62 1.23953205932e-08
L25 139 63 1.07976902515e-08
L26 140 64 1.74396071909e-08
L27 141 65 1.66642462212e-08
L28 142 66 1.48867696727e-08
L29 143 67 1.3105220274e-08
L30 144 68 1.12726810964e-08
L31 145 69 1.19558132861e-08
L32 146 70 1.3165751759e-08
L33 147 71 1.4582803909e-08
L34 148 72 1.61059562721e-08
L35 149 73 1.4712609604e-08
L36 150 74 1.42109542904e-08
L37 151 75 1.38643785983e-08
L38 152 76 1.3712711645e-08
K1_2 L1 L2 0.970037
K1_3 L1 L3 0.93736
K1_4 L1 L4 0.90256
K1_5 L1 L5 0.138112
K1_6 L1 L6 0.124334
K1_7 L1 L7 0.122027
K1_8 L1 L8 0.15667
K1_9 L1 L9 0.140474
K1_10 L1 L10 0.173734
K1_11 L1 L11 0.152738
K1_12 L1 L12 0.177684
K1_13 L1 L13 0.158862
K1_14 L1 L14 0.106751
K1_15 L1 L15 0.121913
K1_16 L1 L16 0.132589
K1_17 L1 L17 0.138453
K1_18 L1 L18 -0.00754008
K1_19 L1 L19 -0.00352049
K1_20 L1 L20 -0.000627933
K1_21 L1 L21 0.00139349
K1_22 L1 L22 0.00288734
K1_23 L1 L23 0.0129383
K1_24 L1 L24 0.0226978
K1_25 L1 L25 0.0310757
K1_26 L1 L26 -0.0122015
K1_27 L1 L27 -0.00482436
K1_28 L1 L28 0.00433152
K1_29 L1 L29 0.0135844
K1_30 L1 L30 0.0218794
K1_31 L1 L31 0.0431703
K1_32 L1 L32 0.006811
K1_33 L1 L33 -0.0325441
K1_34 L1 L34 -0.0738329
K1_35 L1 L35 -0.019496
K1_36 L1 L36 -0.00476307
K1_37 L1 L37 0.00766252
K1_38 L1 L38 0.0167034
K2_3 L2 L3 0.967674
K2_4 L2 L4 0.932032
K2_5 L2 L5 0.139118
K2_6 L2 L6 0.129873
K2_7 L2 L7 0.123967
K2_8 L2 L8 0.159553
K2_9 L2 L9 0.140469
K2_10 L2 L10 0.168983
K2_11 L2 L11 0.148671
K2_12 L2 L12 0.167069
K2_13 L2 L13 0.150986
K2_14 L2 L14 0.107963
K2_15 L2 L15 0.121624
K2_16 L2 L16 0.12917
K2_17 L2 L17 0.132138
K2_18 L2 L18 -0.00636667
K2_19 L2 L19 -0.00234224
K2_20 L2 L20 -0.000119207
K2_21 L2 L21 0.000866692
K2_22 L2 L22 0.0069452
K2_23 L2 L23 0.0161066
K2_24 L2 L24 0.0243292
K2_25 L2 L25 0.0311407
K2_26 L2 L26 -0.00746972
K2_27 L2 L27 -0.000177661
K2_28 L2 L28 0.00834461
K2_29 L2 L29 0.0163779
K2_30 L2 L30 0.023298
K2_31 L2 L31 0.0396481
K2_32 L2 L32 0.0280231
K2_33 L2 L33 -0.00874526
K2_34 L2 L34 -0.0519646
K2_35 L2 L35 -0.0092446
K2_36 L2 L36 0.00428023
K2_37 L2 L37 0.0142129
K2_38 L2 L38 0.0205647
K3_4 L3 L4 0.964623
K3_5 L3 L5 0.138776
K3_6 L3 L6 0.136352
K3_7 L3 L7 0.125104
K3_8 L3 L8 0.157646
K3_9 L3 L9 0.137539
K3_10 L3 L10 0.158849
K3_11 L3 L11 0.14133
K3_12 L3 L12 0.155042
K3_13 L3 L13 0.141521
K3_14 L3 L14 0.108304
K3_15 L3 L15 0.118938
K3_16 L3 L16 0.1231
K3_17 L3 L17 0.124361
K3_18 L3 L18 -0.00469999
K3_19 L3 L19 -0.00129928
K3_20 L3 L20 -4.3494e-05
K3_21 L3 L21 0.000292465
K3_22 L3 L22 0.0115871
K3_23 L3 L23 0.0193887
K3_24 L3 L24 0.0259387
K3_25 L3 L25 0.0315017
K3_26 L3 L26 -0.00210803
K3_27 L3 L27 0.00492301
K3_28 L3 L28 0.0124214
K3_29 L3 L29 0.0190221
K3_30 L3 L30 0.0247251
K3_31 L3 L31 0.0410647
K3_32 L3 L32 0.0345745
K3_33 L3 L33 0.021428
K3_34 L3 L34 -0.0198779
K3_35 L3 L35 0.00699235
K3_36 L3 L36 0.0183126
K3_37 L3 L37 0.0254703
K3_38 L3 L38 0.0299557
K4_5 L4 L5 0.136464
K4_6 L4 L6 0.139302
K4_7 L4 L7 0.123799
K4_8 L4 L8 0.148812
K4_9 L4 L9 0.131042
K4_10 L4 L10 0.147044
K4_11 L4 L11 0.132303
K4_12 L4 L12 0.142983
K4_13 L4 L13 0.13146
K4_14 L4 L14 0.106568
K4_15 L4 L15 0.113384
K4_16 L4 L16 0.115554
K4_17 L4 L17 0.115872
K4_18 L4 L18 -0.00292462
K4_19 L4 L19 -0.000682912
K4_20 L4 L20 -0.000116916
K4_21 L4 L21 -7.39697e-05
K4_22 L4 L22 0.0161853
K4_23 L4 L23 0.02247
K4_24 L4 L24 0.0276934
K4_25 L4 L25 0.0324127
K4_26 L4 L26 0.00343736
K4_27 L4 L27 0.0100255
K4_28 L4 L28 0.0162835
K4_29 L4 L29 0.0216273
K4_30 L4 L30 0.026448
K4_31 L4 L31 0.0443239
K4_32 L4 L32 0.0384147
K4_33 L4 L33 0.0302823
K4_34 L4 L34 0.0123291
K4_35 L4 L35 0.0212811
K4_36 L4 L36 0.0298138
K4_37 L4 L37 0.0349402
K4_38 L4 L38 0.0382795
K5_6 L5 L6 0.780599
K5_7 L5 L7 0.709859
K5_8 L5 L8 0.758333
K5_9 L5 L9 0.689239
K5_10 L5 L10 0.727347
K5_11 L5 L11 0.66744
K5_12 L5 L12 0.694387
K5_13 L5 L13 0.645385
K5_14 L5 L14 0.619708
K5_15 L5 L15 0.604216
K5_16 L5 L16 0.588661
K5_17 L5 L17 0.573218
K5_18 L5 L18 -0.013794
K5_19 L5 L19 -0.0051138
K5_20 L5 L20 -0.00296447
K5_21 L5 L21 -0.00250523
K5_22 L5 L22 0.0251024
K5_23 L5 L23 0.0286088
K5_24 L5 L24 0.0316834
K5_25 L5 L25 0.0353131
K5_26 L5 L26 -0.00198194
K5_27 L5 L27 0.0170852
K5_28 L5 L28 0.0220228
K5_29 L5 L29 0.0252251
K5_30 L5 L30 0.0288023
K5_31 L5 L31 0.0346908
K5_32 L5 L32 0.0278258
K5_33 L5 L33 0.0190825
K5_34 L5 L34 0.0072803
K5_35 L5 L35 0.030034
K5_36 L5 L36 0.0390523
K5_37 L5 L37 0.0424386
K5_38 L5 L38 0.044544
K6_7 L6 L7 0.83362
K6_8 L6 L8 0.93621
K6_9 L6 L9 0.819453
K6_10 L6 L10 0.884605
K6_11 L6 L11 0.79654
K6_12 L6 L12 0.839079
K6_13 L6 L13 0.771895
K6_14 L6 L14 0.705152
K6_15 L6 L15 0.707648
K6_16 L6 L16 0.696453
K6_17 L6 L17 0.681315
K6_18 L6 L18 0.01128
K6_19 L6 L19 0.00712404
K6_20 L6 L20 0.00479059
K6_21 L6 L21 0.00407175
K6_22 L6 L22 0.00775326
K6_23 L6 L23 0.0251823
K6_24 L6 L24 0.035519
K6_25 L6 L25 0.0427484
K6_26 L6 L26 -0.0255891
K6_27 L6 L27 -0.00698768
K6_28 L6 L28 0.013407
K6_29 L6 L29 0.0253626
K6_30 L6 L30 0.0333591
K6_31 L6 L31 0.0160038
K6_32 L6 L32 0.0169505
K6_33 L6 L33 0.018663
K6_34 L6 L34 0.0134697
K6_35 L6 L35 -0.0418814
K6_36 L6 L36 -0.024248
K6_37 L6 L37 -0.016697
K6_38 L6 L38 -0.0123804
K7_8 L7 L8 0.803275
K7_9 L7 L9 0.726904
K7_10 L7 L10 0.764932
K7_11 L7 L11 0.697965
K7_12 L7 L12 0.728026
K7_13 L7 L13 0.674329
K7_14 L7 L14 0.855749
K7_15 L7 L15 0.633256
K7_16 L7 L16 0.613561
K7_17 L7 L17 0.597572
K7_18 L7 L18 0.00428231
K7_19 L7 L19 -0.000496013
K7_20 L7 L20 -0.000367087
K7_21 L7 L21 -0.000398171
K7_22 L7 L22 0.0119577
K7_23 L7 L23 0.0236118
K7_24 L7 L24 0.0296102
K7_25 L7 L25 0.0342649
K7_26 L7 L26 -0.0189637
K7_27 L7 L27 -0.00109281
K7_28 L7 L28 0.0144499
K7_29 L7 L29 0.0219597
K7_30 L7 L30 0.0270567
K7_31 L7 L31 0.0250825
K7_32 L7 L32 0.0205663
K7_33 L7 L33 0.0145263
K7_34 L7 L34 0.00419094
K7_35 L7 L35 0.0081251
K7_36 L7 L36 0.0180074
K7_37 L7 L37 0.0216675
K7_38 L7 L38 0.0241174
K8_9 L8 L9 0.871931
K8_10 L8 L10 0.943232
K8_11 L8 L11 0.850207
K8_12 L8 L12 0.894007
K8_13 L8 L13 0.823504
K8_14 L8 L14 0.682033
K8_15 L8 L15 0.753182
K8_16 L8 L16 0.743256
K8_17 L8 L17 0.727179
K8_18 L8 L18 0.00377852
K8_19 L8 L19 0.00501653
K8_20 L8 L20 0.00421793
K8_21 L8 L21 0.00321289
K8_22 L8 L22 -0.00413603
K8_23 L8 L23 0.0189012
K8_24 L8 L24 0.0321366
K8_25 L8 L25 0.0403206
K8_26 L8 L26 -0.0388941
K8_27 L8 L27 -0.0191754
K8_28 L8 L28 0.00526086
K8_29 L8 L29 0.0204715
K8_30 L8 L30 0.029846
K8_31 L8 L31 0.0209902
K8_32 L8 L32 0.0174846
K8_33 L8 L33 0.00478915
K8_34 L8 L34 -0.0202111
K8_35 L8 L35 -0.0482483
K8_36 L8 L36 -0.0162777
K8_37 L8 L37 -0.00436102
K8_38 L8 L38 0.000631025
K9_10 L9 L10 0.837031
K9_11 L9 L11 0.769456
K9_12 L9 L12 0.79705
K9_13 L9 L13 0.739632
K9_14 L9 L14 0.621813
K9_15 L9 L15 0.868359
K9_16 L9 L16 0.676999
K9_17 L9 L17 0.655841
K9_18 L9 L18 -0.0058039
K9_19 L9 L19 0.000903269
K9_20 L9 L20 -0.00194181
K9_21 L9 L21 -0.00152037
K9_22 L9 L22 -0.00392833
K9_23 L9 L23 0.0179733
K9_24 L9 L24 0.027411
K9_25 L9 L25 0.0329751
K9_26 L9 L26 -0.0364166
K9_27 L9 L27 -0.0175157
K9_28 L9 L28 0.0055315
K9_29 L9 L29 0.0179711
K9_30 L9 L30 0.0246223
K9_31 L9 L31 0.0267549
K9_32 L9 L32 0.0184228
K9_33 L9 L33 0.00497401
K9_34 L9 L34 -0.0143047
K9_35 L9 L35 -0.00886952
K9_36 L9 L36 0.0253733
K9_37 L9 L37 0.0315975
K9_38 L9 L38 0.0342861
K10_11 L10 L11 0.900516
K10_12 L10 L12 0.945935
K10_13 L10 L13 0.871875
K10_14 L10 L14 0.651231
K10_15 L10 L15 0.724611
K10_16 L10 L16 0.78683
K10_17 L10 L17 0.769505
K10_18 L10 L18 -0.00106457
K10_19 L10 L19 -0.00130855
K10_20 L10 L20 0.00257992
K10_21 L10 L21 0.0027542
K10_22 L10 L22 -0.0197771
K10_23 L10 L23 0.00654778
K10_24 L10 L24 0.0269077
K10_25 L10 L25 0.0385367
K10_26 L10 L26 -0.0540673
K10_27 L10 L27 -0.0345267
K10_28 L10 L28 -0.00817729
K10_29 L10 L29 0.0124449
K10_30 L10 L30 0.0257496
K10_31 L10 L31 0.0275832
K10_32 L10 L32 0.0087808
K10_33 L10 L33 -0.0182764
K10_34 L10 L34 -0.0445545
K10_35 L10 L35 -0.0516372
K10_36 L10 L36 -0.0153126
K10_37 L10 L37 0.0129117
K10_38 L10 L38 0.0222406
K11_12 L11 L12 0.860308
K11_13 L11 L13 0.802282
K11_14 L11 L14 0.596477
K11_15 L11 L15 0.669259
K11_16 L11 L16 0.87671
K11_17 L11 L17 0.711875
K11_18 L11 L18 -0.00534541
K11_19 L11 L19 -0.00853515
K11_20 L11 L20 -0.000609834
K11_21 L11 L21 -0.0031946
K11_22 L11 L22 -0.0225655
K11_23 L11 L23 0.00295653
K11_24 L11 L24 0.023189
K11_25 L11 L25 0.0324402
K11_26 L11 L26 -0.0541318
K11_27 L11 L27 -0.0357204
K11_28 L11 L28 -0.0106135
K11_29 L11 L29 0.0097903
K11_30 L11 L30 0.0215715
K11_31 L11 L31 0.0290487
K11_32 L11 L32 0.0121629
K11_33 L11 L33 -0.00930879
K11_34 L11 L34 -0.0311694
K11_35 L11 L35 -0.0191004
K11_36 L11 L36 0.0164149
K11_37 L11 L37 0.0471302
K11_38 L11 L38 0.0522496
K12_13 L12 L13 0.923915
K12_14 L12 L14 0.620622
K12_15 L12 L15 0.691277
K12_16 L12 L16 0.753074
K12_17 L12 L17 0.814397
K12_18 L12 L18 -0.0031561
K12_19 L12 L19 -0.00533954
K12_20 L12 L20 -0.00373198
K12_21 L12 L21 0.00168316
K12_22 L12 L22 -0.0335791
K12_23 L12 L23 -0.00708214
K12_24 L12 L24 0.0174151
K12_25 L12 L25 0.0376503
K12_26 L12 L26 -0.067791
K12_27 L12 L27 -0.0490397
K12_28 L12 L28 -0.0230335
K12_29 L12 L29 0.000206869
K12_30 L12 L30 0.0199571
K12_31 L12 L31 0.0265907
K12_32 L12 L32 -0.00333105
K12_33 L12 L33 -0.0313495
K12_34 L12 L34 -0.0564259
K12_35 L12 L35 -0.0438762
K12_36 L12 L36 -0.00790358
K12_37 L12 L37 0.0248258
K12_38 L12 L38 0.0534953
K13_14 L13 L14 0.576034
K13_15 L13 L15 0.642945
K13_16 L13 L16 0.704816
K13_17 L13 L17 0.884083
K13_18 L13 L18 -0.00514509
K13_19 L13 L19 -0.00824098
K13_20 L13 L20 -0.00977699
K13_21 L13 L21 -0.00215163
K13_22 L13 L22 -0.0370798
K13_23 L13 L23 -0.0119354
K13_24 L13 L24 0.0122548
K13_25 L13 L25 0.0329791
K13_26 L13 L26 -0.0685963
K13_27 L13 L27 -0.0509855
K13_28 L13 L28 -0.0264989
K13_29 L13 L29 -0.00381141
K13_30 L13 L30 0.0162576
K13_31 L13 L31 0.0281607
K13_32 L13 L32 0.00369445
K13_33 L13 L33 -0.0202422
K13_34 L13 L34 -0.042551
K13_35 L13 L35 -0.0123318
K13_36 L13 L36 0.0222888
K13_37 L13 L37 0.0545038
K13_38 L13 L38 0.0849571
K14_15 L14 L15 0.547961
K14_16 L14 L16 0.526055
K14_17 L14 L17 0.511368
K14_18 L14 L18 -0.115303
K14_19 L14 L19 -0.0074497
K14_20 L14 L20 -0.00268917
K14_21 L14 L21 -0.00181956
K14_22 L14 L22 0.0133953
K14_23 L14 L23 0.0203328
K14_24 L14 L24 0.024275
K14_25 L14 L25 0.0277337
K14_26 L14 L26 -0.0178823
K14_27 L14 L27 0.00312225
K14_28 L14 L28 0.0136536
K14_29 L14 L29 0.0184181
K14_30 L14 L30 0.0220779
K14_31 L14 L31 0.0239192
K14_32 L14 L32 0.0191755
K14_33 L14 L33 0.0130015
K14_34 L14 L34 0.00333841
K14_35 L14 L35 0.0126797
K14_36 L14 L36 0.023079
K14_37 L14 L37 0.0263943
K14_38 L14 L38 0.0283916
K15_16 L15 L16 0.59432
K15_17 L15 L17 0.571621
K15_18 L15 L18 -0.0211377
K15_19 L15 L19 -0.112503
K15_20 L15 L20 -0.00830095
K15_21 L15 L21 -0.00362575
K15_22 L15 L22 -0.00188478
K15_23 L15 L23 0.0171391
K15_24 L15 L24 0.0226997
K15_25 L15 L25 0.0266157
K15_26 L15 L26 -0.0317861
K15_27 L15 L27 -0.0142668
K15_28 L15 L28 0.00710984
K15_29 L15 L29 0.0157252
K15_30 L15 L30 0.0201798
K15_31 L15 L31 0.0250364
K15_32 L15 L32 0.0172568
K15_33 L15 L33 0.00533241
K15_34 L15 L34 -0.0112806
K15_35 L15 L35 0.000402055
K15_36 L15 L36 0.0271307
K15_37 L15 L37 0.0343952
K15_38 L15 L38 0.0369936
K16_17 L16 L17 0.630701
K16_18 L16 L18 -0.00813642
K16_19 L16 L19 -0.0227781
K16_20 L16 L20 -0.110447
K16_21 L16 L21 -0.00972946
K16_22 L16 L22 -0.0221385
K16_23 L16 L23 0.00136233
K16_24 L16 L24 0.0191767
K16_25 L16 L25 0.0247684
K16_26 L16 L26 -0.0501204
K16_27 L16 L27 -0.0335874
K16_28 L16 L28 -0.0107575
K16_29 L16 L29 0.0087675
K16_30 L16 L30 0.0171848
K16_31 L16 L31 0.0269264
K16_32 L16 L32 0.0122878
K16_33 L16 L33 -0.00606963
K16_34 L16 L34 -0.0248461
K16_35 L16 L35 -0.0080866
K16_36 L16 L36 0.0228636
K16_37 L16 L37 0.0468301
K16_38 L16 L38 0.0531762
K17_18 L17 L18 -0.00621429
K17_19 L17 L19 -0.0106781
K17_20 L17 L20 -0.0238487
K17_21 L17 L21 -0.109989
K17_22 L17 L22 -0.0429948
K17_23 L17 L23 -0.0207529
K17_24 L17 L24 0.00153511
K17_25 L17 L25 0.0200322
K17_26 L17 L26 -0.0677959
K17_27 L17 L27 -0.0521188
K17_28 L17 L28 -0.0304093
K17_29 L17 L29 -0.00955488
K17_30 L17 L30 0.00998879
K17_31 L17 L31 0.0265623
K17_32 L17 L32 0.00587095
K17_33 L17 L33 -0.0146158
K17_34 L17 L34 -0.0340072
K17_35 L17 L35 -0.000672041
K17_36 L17 L36 0.0303199
K17_37 L17 L37 0.0586492
K17_38 L17 L38 0.0825751
K18_19 L18 L19 0.018364
K18_20 L18 L20 0.00503238
K18_21 L18 L21 0.00290319
K18_22 L18 L22 0.00115055
K18_23 L18 L23 3.55839e-05
K18_24 L18 L24 0.00152562
K18_25 L18 L25 0.00209948
K18_26 L18 L26 0.0078735
K18_27 L18 L27 0.00209275
K18_28 L18 L28 -0.000666932
K18_29 L18 L29 0.0010789
K18_30 L18 L30 0.00190822
K18_31 L18 L31 -0.00396486
K18_32 L18 L32 -0.00174985
K18_33 L18 L33 0.00080015
K18_34 L18 L34 0.00305024
K18_35 L18 L35 -0.00247983
K18_36 L18 L36 -0.01236
K18_37 L18 L37 -0.0139724
K18_38 L18 L38 -0.0142729
K19_20 L19 L20 0.0186651
K19_21 L19 L21 0.00546108
K19_22 L19 L22 0.0100611
K19_23 L19 L23 0.0032237
K19_24 L19 L24 0.00154314
K19_25 L19 L25 0.00260731
K19_26 L19 L26 0.0100038
K19_27 L19 L27 0.00875163
K19_28 L19 L28 0.00461413
K19_29 L19 L29 0.00093764
K19_30 L19 L30 0.00224786
K19_31 L19 L31 -0.00345127
K19_32 L19 L32 -0.00135286
K19_33 L19 L33 0.000150102
K19_34 L19 L34 0.000812341
K19_35 L19 L35 -0.00416473
K19_36 L19 L36 -0.00422605
K19_37 L19 L37 -0.014261
K19_38 L19 L38 -0.0160491
K20_21 L20 L21 0.0200064
K20_22 L20 L22 0.015979
K20_23 L20 L23 0.0145528
K20_24 L20 L24 0.00717083
K20_25 L20 L25 0.00493259
K20_26 L20 L26 0.0140842
K20_27 L20 L27 0.0137741
K20_28 L20 L28 0.0127608
K20_29 L20 L29 0.00810448
K20_30 L20 L30 0.00374733
K20_31 L20 L31 -0.00286489
K20_32 L20 L32 -0.00192188
K20_33 L20 L33 -0.00179125
K20_34 L20 L34 -0.00187392
K20_35 L20 L35 -0.00693624
K20_36 L20 L36 -0.0074238
K20_37 L20 L37 -0.00766263
K20_38 L20 L38 -0.0179188
K21_22 L21 L22 0.0225105
K21_23 L21 L23 0.0225789
K21_24 L21 L24 0.0208196
K21_25 L21 L25 0.011704
K21_26 L21 L26 0.0214739
K21_27 L21 L27 0.021518
K21_28 L21 L28 0.021752
K21_29 L21 L29 0.0205519
K21_30 L21 L30 0.0148169
K21_31 L21 L31 -0.00327028
K21_32 L21 L32 -0.00397316
K21_33 L21 L33 -0.00456616
K21_34 L21 L34 -0.00479909
K21_35 L21 L35 -0.014872
K21_36 L21 L36 -0.0158071
K21_37 L21 L37 -0.0166682
K21_38 L21 L38 -0.017109
K22_23 L22 L23 0.947468
K22_24 L22 L24 0.892131
K22_25 L22 L25 0.832903
K22_26 L22 L26 0.307342
K22_27 L22 L27 0.316125
K22_28 L22 L28 0.312762
K22_29 L22 L29 0.304423
K22_30 L22 L30 0.297926
K22_31 L22 L31 0.0149462
K22_32 L22 L32 0.0197734
K22_33 L22 L33 0.0242587
K22_34 L22 L34 0.0276096
K22_35 L22 L35 0.0360182
K22_36 L22 L36 0.0197613
K22_37 L22 L37 -0.000626597
K22_38 L22 L38 -0.0187784
K23_24 L23 L24 0.941488
K23_25 L23 L25 0.878928
K23_26 L23 L26 0.297724
K23_27 L23 L27 0.306163
K23_28 L23 L28 0.323587
K23_29 L23 L29 0.320402
K23_30 L23 L30 0.313485
K23_31 L23 L31 0.0169488
K23_32 L23 L32 0.0200375
K23_33 L23 L33 0.0223855
K23_34 L23 L34 0.0236496
K23_35 L23 L35 0.0247929
K23_36 L23 L36 0.0221915
K23_37 L23 L37 0.00530712
K23_38 L23 L38 -0.0129945
K24_25 L24 L25 0.933592
K24_26 L24 L26 0.287946
K24_27 L24 L27 0.296147
K24_28 L24 L28 0.313009
K24_29 L24 L29 0.332775
K24_30 L24 L30 0.331258
K24_31 L24 L31 0.0195608
K24_32 L24 L32 0.0199218
K24_33 L24 L33 0.0197907
K24_34 L24 L34 0.0193833
K24_35 L24 L35 0.0146186
K24_36 L24 L36 0.0142627
K24_37 L24 L37 0.012081
K24_38 L24 L38 -0.00234193
K25_26 L25 L26 0.27585
K25_27 L25 L27 0.283916
K25_28 L25 L28 0.300161
K25_29 L25 L29 0.31916
K25_30 L25 L30 0.34345
K25_31 L25 L31 0.0220884
K25_32 L25 L32 0.0197297
K25_33 L25 L33 0.0177965
K25_34 L25 L34 0.0163137
K25_35 L25 L35 0.00808453
K25_36 L25 L36 0.00822625
K25_37 L25 L37 0.00872154
K25_38 L25 L38 0.0103187
K26_27 L26 L27 0.976245
K26_28 L26 L28 0.924352
K26_29 L26 L29 0.86907
K26_30 L26 L30 0.809842
K26_31 L26 L31 0.0118477
K26_32 L26 L32 0.0184304
K26_33 L26 L33 0.0244963
K26_34 L26 L34 0.0296176
K26_35 L26 L35 0.0272191
K26_36 L26 L36 0.0107869
K26_37 L26 L37 -0.00652292
K26_38 L26 L38 -0.0228897
K27_28 L27 L28 0.946901
K27_29 L27 L29 0.890245
K27_30 L27 L30 0.829755
K27_31 L27 L31 0.0142343
K27_32 L27 L32 0.02024
K27_33 L27 L33 0.0255334
K27_34 L27 L34 0.0296906
K27_35 L27 L35 0.0289189
K27_36 L27 L36 0.0143427
K27_37 L27 L37 -0.00287663
K27_38 L27 L38 -0.0194286
K28_29 L28 L29 0.940813
K28_30 L28 L30 0.87684
K28_31 L28 L31 0.0159064
K28_32 L28 L32 0.0205818
K28_33 L28 L33 0.0242029
K28_34 L28 L34 0.0266012
K28_35 L28 L35 0.0227821
K28_36 L28 L36 0.0168439
K28_37 L28 L37 0.00146547
K28_38 L28 L38 -0.0152402
K29_30 L29 L30 0.932595
K29_31 L29 L31 0.0183249
K29_32 L29 L32 0.0207779
K29_33 L29 L33 0.0222327
K29_34 L29 L34 0.0229834
K29_35 L29 L35 0.0161368
K29_36 L29 L36 0.0143362
K29_37 L29 L37 0.00817186
K29_38 L29 L38 -0.00654716
K30_31 L30 L31 0.0209878
K30_32 L30 L32 0.0210105
K30_33 L30 L33 0.0206576
K30_34 L30 L34 0.0202468
K30_35 L30 L35 0.0123149
K30_36 L30 L36 0.0114746
K30_37 L30 L37 0.00980212
K30_38 L30 L38 0.00498788
K31_32 L31 L32 0.788887
K31_33 L31 L33 0.743809
K31_34 L31 L34 0.707941
K31_35 L31 L35 0.720271
K31_36 L31 L36 0.734727
K31_37 L31 L37 0.746217
K31_38 L31 L38 0.751557
K32_33 L32 L33 0.808708
K32_34 L32 L34 0.767476
K32_35 L32 L35 0.704436
K32_36 L32 L36 0.716019
K32_37 L32 L37 0.722787
K32_38 L32 L38 0.723495
K33_34 L33 L34 0.826514
K33_35 L33 L35 0.687652
K33_36 L33 L36 0.695122
K33_37 L33 L37 0.697387
K33_38 L33 L38 0.695531
K34_35 L34 L35 0.668875
K34_36 L34 L36 0.671929
K34_37 L34 L37 0.671465
K34_38 L34 L38 0.668299
K35_36 L35 L36 0.975684
K35_37 L35 L37 0.950726
K35_38 L35 L38 0.925053
K36_37 L36 L37 0.974921
K36_38 L36 L38 0.949033
K37_38 L37 L38 0.974221
.ends Quadraat_0004__7_0_6_0_5_0_4_series
.ends Quadraat_0004__7_0_6_0_5_0_4
