* BEGIN ANSOFT HEADER
* node 1    DCPLUS:DCPLUS_LLOAD
* node 2    DCPLUS:DCPLUS_SCAP
* node 3    DCPLUS:DCPLUS_TOPFET
* node 4    GDOUT:Source_GDOUT
* node 5    GND:DCMIN_ISHUNT
* node 6    GND:DCMIN_SCAP
* node 7    GNDM:Kelvin_Source
* node 8    GNDM_2:ISHUNT_SOURCE
* node 9    LOWGATE:Source_TG
* node 10   MIDPOINT:L_SOURCE
* node 11   MIDPOINT:LOWDRN_SOURCE
* node 12   MIDPOINT:VMEAS_SOURCE
* node 13   Vgdl_:GDH_Source
* node 14   DCPLUS:DCPLUS_BIGCAP
* node 15   GDOUT:Sink_GDOUT
* node 16   GND:DCMIN_BIGCAP
* node 17   GNDM:BypassCapGnd
* node 18   GNDM_2:ISHUNT_SINK
* node 19   LOWGATE:Sink_TG
* node 20   MIDPOINT:TOPSRC_SINK
* node 21   Vgdl_:GDH_SINK
*  Project: DPT_PCB3_1
*   Design: Q3DModel1
*   Format: Ansys Nexxim
*   Topckt: DPT_PCB3_1_800kHz
*     Left: 1 2 3 4 5 6 7 8 9 10 11 12 13
*    Right: 14 15 16 17 18 19 20 21
*  Creator: Ansys Electronics Desktop 2021.2.0
*     Date: Fri May 27 00:27:58 2022
* END ANSOFT HEADER

.subckt DPT_PCB3_1_800kHz 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21
XZhalf1 1 2 3 4 5 6 7 8 9 10 11 12 13 27 28 29 30 31 32 33 34 35 36 37 38 39
+ DPT_PCB3_1_800kHz_half
XY1 27 28 29 30 31 32 33 34 35 36 37 38 39 DPT_PCB3_1_800kHz_parlel
XZhalf2 27 28 29 30 31 32 33 34 35 36 37 38 39 14 14 14 15 16 16 17 18 19 20 20
+ 20 21 DPT_PCB3_1_800kHz_half

.subckt DPT_PCB3_1_800kHz_half 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19
+ 20 21 22 23 24 25 26
V1 1 27 dc 0.0
V2 2 28 dc 0.0
V3 3 29 dc 0.0
V4 4 30 dc 0.0
V5 5 31 dc 0.0
V6 6 32 dc 0.0
V7 7 33 dc 0.0
V8 8 34 dc 0.0
V9 9 35 dc 0.0
V10 10 36 dc 0.0
V11 11 37 dc 0.0
V12 12 38 dc 0.0
V13 13 39 dc 0.0
R1 27 40 0.00381516713581
R2 28 41 0.00630583766073
R3 29 42 0.00445334336406
R4 30 43 0.00373264980579
R5 31 44 0.0037554272218
R6 32 45 0.0057898557693
R7 33 46 0.00208700264078
R8 34 47 0.00435469442072
R9 35 48 0.00464951277194
R10 36 49 0.0132888247248
R11 37 50 0.0098354311237
R12 38 51 0.0172727463706
R13 39 52 0.00385491373189
F1_2 40 27 V2 0.520876
F1_3 40 27 V3 0.965508
F1_4 40 27 V4 -0.00716321
F1_5 40 27 V5 0.044446
F1_6 40 27 V6 0.0262643
F1_7 40 27 V7 -0.0233758
F1_8 40 27 V8 0.0192946
F1_9 40 27 V9 -0.00692268
F1_10 40 27 V10 0.0812155
F1_11 40 27 V11 -0.0193915
F1_12 40 27 V12 0.00765571
F1_13 40 27 V13 0.00245997
F2_1 41 28 V1 0.315141
F2_3 41 28 V3 0.3145
F2_4 41 28 V4 -0.00216103
F2_5 41 28 V5 0.0122629
F2_6 41 28 V6 0.00272893
F2_7 41 28 V7 -0.00541214
F2_8 41 28 V8 0.00990959
F2_9 41 28 V9 -0.00174563
F2_10 41 28 V10 0.013392
F2_11 41 28 V11 -0.00538945
F2_12 41 28 V12 0.00488996
F2_13 41 28 V13 6.58554e-05
F3_1 42 29 V1 0.827148
F3_2 42 29 V2 0.445325
F3_4 42 29 V4 -0.00708163
F3_5 42 29 V5 0.0430309
F3_6 42 29 V6 0.0235543
F3_7 42 29 V7 -0.00799889
F3_8 42 29 V8 0.014488
F3_9 42 29 V9 -0.0054643
F3_10 42 29 V10 0.0291755
F3_11 42 29 V11 0.0360526
F3_12 42 29 V12 0.0602551
F3_13 42 29 V13 0.0016854
F4_1 43 30 V1 -0.00732157
F4_2 43 30 V2 -0.00365079
F4_3 43 30 V3 -0.00844894
F4_5 43 30 V5 -0.00735493
F4_6 43 30 V6 -0.00621239
F4_7 43 30 V7 0.0194342
F4_8 43 30 V8 -0.00515469
F4_9 43 30 V9 0.0116512
F4_10 43 30 V10 -0.00377572
F4_11 43 30 V11 -0.0041902
F4_12 43 30 V12 -0.0125328
F4_13 43 30 V13 -0.0262322
F5_1 44 31 V1 0.045153
F5_2 44 31 V2 0.0205909
F5_3 44 31 V3 0.0510279
F5_4 44 31 V4 -0.00731032
F5_6 44 31 V6 0.99505
F5_7 44 31 V7 -0.0140336
F5_8 44 31 V8 0.0150649
F5_9 44 31 V9 -0.00566996
F5_10 44 31 V10 0.0260809
F5_11 44 31 V11 -0.00930359
F5_12 44 31 V12 0.00635412
F5_13 44 31 V13 0.00228831
F6_1 45 32 V1 0.0173066
F6_2 45 32 V2 0.00297213
F6_3 45 32 V3 0.0181171
F6_4 45 32 V4 -0.00400505
F6_5 45 32 V5 0.645411
F6_7 45 32 V7 -0.00714339
F6_8 45 32 V8 0.00691786
F6_9 45 32 V9 -0.00277097
F6_10 45 32 V10 0.0119818
F6_11 45 32 V11 -0.0101545
F6_12 45 32 V12 0.000963965
F6_13 45 32 V13 0.000654648
F7_1 46 33 V1 -0.0427325
F7_2 46 33 V2 -0.0163527
F7_3 46 33 V3 -0.0170684
F7_4 46 33 V4 0.0347585
F7_5 46 33 V5 -0.0252526
F7_6 46 33 V6 -0.0198175
F7_8 46 33 V8 -0.0193199
F7_9 46 33 V9 0.0460094
F7_10 46 33 V10 -0.0232242
F7_11 46 33 V11 -0.0758908
F7_12 46 33 V12 -0.153085
F7_13 46 33 V13 -0.0520915
F8_1 47 34 V1 0.0169041
F8_2 47 34 V2 0.0143496
F8_3 47 34 V3 0.0148162
F8_4 47 34 V4 -0.00441837
F8_5 47 34 V5 0.0129918
F8_6 47 34 V6 0.00919775
F8_7 47 34 V7 -0.00925912
F8_9 47 34 V9 -0.00751556
F8_10 47 34 V10 0.0219934
F8_11 47 34 V11 0.0183315
F8_12 47 34 V12 0.0525452
F8_13 47 34 V13 0.00256465
F9_1 48 35 V1 -0.00568042
F9_2 48 35 V2 -0.00236749
F9_3 48 35 V3 -0.00523376
F9_4 48 35 V4 0.00935366
F9_5 48 35 V5 -0.00457965
F9_6 48 35 V6 -0.00345058
F9_7 48 35 V7 0.020652
F9_8 48 35 V8 -0.00703901
F9_10 48 35 V10 -0.00189503
F9_11 48 35 V11 -0.0159624
F9_12 48 35 V12 -0.0229492
F9_13 48 35 V13 -0.00811278
F10_1 49 36 V1 0.0233166
F10_2 49 36 V2 0.00635482
F10_3 49 36 V3 0.00977727
F10_4 49 36 V4 -0.00106055
F10_5 49 36 V5 0.00737047
F10_6 49 36 V6 0.00522041
F10_7 49 36 V7 -0.00364735
F10_8 49 36 V8 0.00720715
F10_9 49 36 V9 -0.000663035
F10_11 49 36 V11 0.0434243
F10_12 49 36 V12 0.0509842
F10_13 49 36 V13 -0.000873577
F11_1 50 37 V1 -0.00752196
F11_2 50 37 V2 -0.00345536
F11_3 50 37 V3 0.0163241
F11_4 50 37 V4 -0.00159023
F11_5 50 37 V5 -0.00355236
F11_6 50 37 V6 -0.00597769
F11_7 50 37 V7 -0.0161034
F11_8 50 37 V8 0.00811639
F11_9 50 37 V9 -0.00754592
F11_10 50 37 V10 0.0586714
F11_12 50 37 V12 0.989122
F11_13 50 37 V13 0.00524892
F12_1 51 38 V1 0.00169098
F12_2 51 38 V2 0.0017852
F12_3 51 38 V3 0.0155353
F12_4 51 38 V4 -0.00270834
F12_5 51 38 V5 0.00138151
F12_6 51 38 V6 0.000323123
F12_7 51 38 V7 -0.0184967
F12_8 51 38 V8 0.0132474
F12_9 51 38 V9 -0.00617751
F12_10 51 38 V10 0.0392248
F12_11 51 38 V11 0.563225
F12_13 51 38 V13 0.00405379
F13_1 52 39 V1 0.0024346
F13_2 52 39 V2 0.000107726
F13_3 52 39 V3 0.00194704
F13_4 52 39 V4 -0.0254002
F13_5 52 39 V5 0.00222926
F13_6 52 39 V6 0.000983243
F13_7 52 39 V7 -0.0282017
F13_8 52 39 V8 0.00289716
F13_9 52 39 V9 -0.00978504
F13_10 52 39 V10 -0.00301143
F13_11 52 39 V11 0.0133921
F13_12 52 39 V12 0.0181638
L1 40 14 1.33468306618e-08
L2 41 15 6.56906069955e-09
L3 42 16 1.44986646669e-08
L4 43 17 1.11831507759e-09
L5 44 18 8.00061715858e-09
L6 45 19 8.38185844268e-09
L7 46 20 1.71983847127e-09
L8 47 21 3.3257344411e-09
L9 48 22 1.70653836206e-09
L10 49 23 1.09135164766e-08
L11 50 24 7.08825700825e-09
L12 51 25 1.17906826613e-08
L13 52 26 1.19335663402e-09
K1_2 L1 L2 0.575098
K1_3 L1 L3 0.927058
K1_4 L1 L4 -0.0150628
K1_5 L1 L5 0.0708412
K1_6 L1 L6 0.0585372
K1_7 L1 L7 -0.0297254
K1_8 L1 L8 0.0211151
K1_9 L1 L9 -0.00988022
K1_10 L1 L10 0.073796
K1_11 L1 L11 -0.00711991
K1_12 L1 L12 0.0161212
K1_13 L1 L13 0.00415304
K2_3 L2 L3 0.54956
K2_4 L2 L4 -0.00838748
K2_5 L2 L5 0.0617322
K2_6 L2 L6 0.0515349
K2_7 L2 L7 -0.0154873
K2_8 L2 L8 0.0119135
K2_9 L2 L9 -0.00487085
K2_10 L2 L10 0.0249371
K2_11 L2 L11 -0.00500029
K2_12 L2 L12 0.00712059
K2_13 L2 L13 0.00169707
K3_4 L3 L4 -0.0159318
K3_5 L3 L5 0.071946
K3_6 L3 L6 0.059751
K3_7 L3 L7 -0.0330983
K3_8 L3 L8 0.0228701
K3_9 L3 L9 -0.0140586
K3_10 L3 L10 0.0133976
K3_11 L3 L11 0.0231224
K3_12 L3 L12 0.0395108
K3_13 L3 L13 0.00745782
K4_5 L4 L5 -0.0176032
K4_6 L4 L6 -0.0156297
K4_7 L4 L7 0.0919081
K4_8 L4 L8 -0.0133582
K4_9 L4 L9 0.0237168
K4_10 L4 L10 -0.00878848
K4_11 L4 L11 -4.87041e-05
K4_12 L4 L12 -0.0293612
K4_13 L4 L13 -0.178112
K5_6 L5 L6 0.946286
K5_7 L5 L7 -0.0341227
K5_8 L5 L8 0.0194798
K5_9 L5 L9 -0.0143541
K5_10 L5 L10 0.0132411
K5_11 L5 L11 0.00155494
K5_12 L5 L12 0.0177131
K5_13 L5 L13 0.00837739
K6_7 L6 L7 -0.0298165
K6_8 L6 L8 0.0152032
K6_9 L6 L9 -0.0125753
K6_10 L6 L10 0.0107077
K6_11 L6 L11 0.0012724
K6_12 L6 L12 0.0153519
K6_13 L6 L13 0.0075793
K7_8 L7 L8 -0.0440951
K7_9 L7 L9 0.341218
K7_10 L7 L10 -0.012382
K7_11 L7 L11 -0.022252
K7_12 L7 L12 -0.144699
K7_13 L7 L13 -0.0704012
K8_9 L8 L9 -0.0270874
K8_10 L8 L10 0.00969701
K8_11 L8 L11 0.0116025
K8_12 L8 L12 0.0391514
K8_13 L8 L13 0.00736605
K9_10 L9 L10 -0.0014249
K9_11 L9 L11 -0.0167204
K9_12 L9 L12 -0.0633161
K9_13 L9 L13 -0.0381987
K10_11 L10 L11 -0.0102429
K10_12 L10 L12 0.0109177
K10_13 L10 L13 -0.00164266
K11_12 L11 L12 0.760154
K11_13 L11 L13 0.0118526
K12_13 L12 L13 0.0245961
.ends DPT_PCB3_1_800kHz_half

.subckt DPT_PCB3_1_800kHz_parlel 1 2 3 4 5 6 7 8 9 10 11 12 13
RG1_4 1 4 -1.98350110422e+12
RG1_5 1 5 108575247.199
RG1_6 1 6 108575247.199
RG1_7 1 7 61006775825.9
RG1_8 1 8 1466265290.65
RG1_9 1 9 311003448140
RG1_10 1 10 1049784358.77
RG1_11 1 11 1049784358.77
RG1_12 1 12 1049784358.77
RG1_13 1 13 -188399965979
RG2_4 2 4 -1.98350110422e+12
RG2_5 2 5 108575247.199
RG2_6 2 6 108575247.199
RG2_7 2 7 61006775825.9
RG2_8 2 8 1466265290.65
RG2_9 2 9 311003448140
RG2_10 2 10 1049784358.77
RG2_11 2 11 1049784358.77
RG2_12 2 12 1049784358.77
RG2_13 2 13 -188399965979
RG3_4 3 4 -1.98350110422e+12
RG3_5 3 5 108575247.199
RG3_6 3 6 108575247.199
RG3_7 3 7 61006775825.9
RG3_8 3 8 1466265290.65
RG3_9 3 9 311003448140
RG3_10 3 10 1049784358.77
RG3_11 3 11 1049784358.77
RG3_12 3 12 1049784358.77
RG3_13 3 13 -188399965979
R4_0 4 0 28328705.4553
RG4_5 4 5 3.23224702611e+12
RG4_6 4 6 3.23224702611e+12
RG4_7 4 7 286576194.166
RG4_8 4 8 -1.18367652795e+12
RG4_9 4 9 -245544099753
RG4_10 4 10 -967418316797
RG4_11 4 11 -967418316797
RG4_12 4 12 -967418316797
RG4_13 4 13 77316092.8419
R5_0 5 0 1740542961.7
RG5_7 5 7 1207286403.33
RG5_8 5 8 66982279.2231
RG5_9 5 9 -53078935390
RG5_10 5 10 44820735354.5
RG5_11 5 11 44820735354.5
RG5_12 5 12 44820735354.5
RG5_13 5 13 104706073276
R6_0 6 0 1740542961.7
RG6_7 6 7 1207286403.33
RG6_8 6 8 66982279.2231
RG6_9 6 9 -53078935390
RG6_10 6 10 44820735354.5
RG6_11 6 11 44820735354.5
RG6_12 6 12 44820735354.5
RG6_13 6 13 104706073276
R7_0 7 0 3189714.61286
RG7_8 7 8 44139048.436
RG7_9 7 9 5114925.35817
RG7_10 7 10 110511852.142
RG7_11 7 11 110511852.142
RG7_12 7 12 110511852.142
RG7_13 7 13 7724579.85831
R8_0 8 0 754357553.773
RG8_9 8 9 5.58283056e+12
RG8_10 8 10 730388308.019
RG8_11 8 11 730388308.019
RG8_12 8 12 730388308.019
RG8_13 8 13 -202932013606
RG9_10 9 10 -145085276597
RG9_11 9 11 -145085276597
RG9_12 9 12 -145085276597
RG9_13 9 13 -206506194866
R10_0 10 0 180291762.569
RG10_13 10 13 255471858425
R11_0 11 0 180291762.569
RG11_13 11 13 255471858425
R12_0 12 0 180291762.569
RG12_13 12 13 255471858425
R13_0 13 0 216828764.481
C1_0 1 0 5.14712751185e-13
C1_4 1 4 6.28947727255e-17
C1_5 1 5 4.69657696703e-13
C1_6 1 6 4.69657696703e-13
C1_7 1 7 1.25321953336e-13
C1_8 1 8 6.60420159676e-14
C1_9 1 9 7.39212429332e-16
C1_10 1 10 4.17893138593e-14
C1_11 1 11 4.17893138593e-14
C1_12 1 12 4.17893138593e-14
C1_13 1 13 1.11026862323e-15
C2_0 2 0 5.14712751185e-13
C2_4 2 4 6.28947727255e-17
C2_5 2 5 4.69657696703e-13
C2_6 2 6 4.69657696703e-13
C2_7 2 7 1.25321953336e-13
C2_8 2 8 6.60420159676e-14
C2_9 2 9 7.39212429332e-16
C2_10 2 10 4.17893138593e-14
C2_11 2 11 4.17893138593e-14
C2_12 2 12 4.17893138593e-14
C2_13 2 13 1.11026862323e-15
C3_0 3 0 5.14712751185e-13
C3_4 3 4 6.28947727255e-17
C3_5 3 5 4.69657696703e-13
C3_6 3 6 4.69657696703e-13
C3_7 3 7 1.25321953336e-13
C3_8 3 8 6.60420159676e-14
C3_9 3 9 7.39212429332e-16
C3_10 3 10 4.17893138593e-14
C3_11 3 11 4.17893138593e-14
C3_12 3 12 4.17893138593e-14
C3_13 3 13 1.11026862323e-15
C4_0 4 0 4.53704708796e-13
C4_5 4 5 2.00013463255e-16
C4_6 4 6 2.00013463255e-16
C4_7 4 7 7.38047047522e-14
C4_8 4 8 2.34285898609e-16
C4_9 4 9 1.63342773226e-16
C4_10 4 10 4.99653088882e-17
C4_11 4 11 4.99653088882e-17
C4_12 4 12 4.99653088882e-17
C4_13 4 13 1.77927388535e-13
C5_0 5 0 7.30927844047e-13
C5_7 5 7 2.75959105827e-13
C5_8 5 8 5.52363114015e-13
C5_9 5 9 2.08021148626e-15
C5_10 5 10 8.98078766663e-15
C5_11 5 11 8.98078766663e-15
C5_12 5 12 8.98078766663e-15
C5_13 5 13 2.41416714297e-15
C6_0 6 0 7.30927844047e-13
C6_7 6 7 2.75959105827e-13
C6_8 6 8 5.52363114015e-13
C6_9 6 9 2.08021148626e-15
C6_10 6 10 8.98078766663e-15
C6_11 6 11 8.98078766663e-15
C6_12 6 12 8.98078766663e-15
C6_13 6 13 2.41416714297e-15
C7_0 7 0 6.01517021414e-12
C7_8 7 8 7.56655046778e-13
C7_9 7 9 2.66402134727e-12
C7_10 7 10 3.11587561308e-13
C7_11 7 11 3.11587561308e-13
C7_12 7 12 3.11587561308e-13
C7_13 7 13 2.46623901856e-12
C8_0 8 0 1.3410363457e-13
C8_9 8 9 1.08975701455e-14
C8_10 8 10 5.22320901808e-14
C8_11 8 11 5.22320901808e-14
C8_12 8 12 5.22320901808e-14
C8_13 8 13 1.92931468429e-15
C9_10 9 10 1.42277168824e-15
C9_11 9 11 1.42277168824e-15
C9_12 9 12 1.42277168824e-15
C9_13 9 13 7.22422118735e-16
C10_0 10 0 1.65565373774e-13
C10_13 10 13 9.91456088168e-16
C11_0 11 0 1.65565373774e-13
C11_13 11 13 9.91456088168e-16
C12_0 12 0 1.65565373774e-13
C12_13 12 13 9.91456088168e-16
C13_0 13 0 1.34765793868e-13
.ends DPT_PCB3_1_800kHz_parlel

.ends DPT_PCB3_1_800kHz
