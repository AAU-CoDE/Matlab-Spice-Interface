* BEGIN ANSOFT HEADER
* node 1    DCPLUS:DCPLUS_LLOAD
* node 2    DCPLUS:DCPLUS_SCAP
* node 3    DCPLUS:DCPLUS_TOPFET
* node 4    GDOUT:Source_GDOUT
* node 5    GND:DCMIN_ISHUNT
* node 6    GND:DCMIN_SCAP
* node 7    GNDM:Kelvin_Source
* node 8    GNDM_2:ISHUNT_SOURCE
* node 9    LOWGATE:Source_TG
* node 10   MIDPOINT:L_SOURCE
* node 11   MIDPOINT:LOWDRN_SOURCE
* node 12   MIDPOINT:VMEAS_SOURCE
* node 13   Vgdl_:GDH_Source
* node 14   DCPLUS:DCPLUS_BIGCAP
* node 15   GDOUT:Sink_GDOUT
* node 16   GND:DCMIN_BIGCAP
* node 17   GNDM:BypassCapGnd
* node 18   GNDM_2:ISHUNT_SINK
* node 19   LOWGATE:Sink_TG
* node 20   MIDPOINT:TOPSRC_SINK
* node 21   Vgdl_:GDH_SINK
*  Project: DPT_PCB2
*   Design: Q3DModel1
*   Format: ANSYS Nexxim
*   Topckt: DPT_PCB3_1MHz
*     Left: 1 2 3 4 5 6 7 8 9 10 11 12 13
*    Right: 14 15 16 17 18 19 20 21
*  Creator: Ansoft Electronics Desktop 2021.1.0
*     Date: Sun Mar 06 15:48:33 2022
* END ANSOFT HEADER

.subckt DPT_PCB3_1MHz 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21
XZhalf1 1 2 3 4 5 6 7 8 9 10 11 12 13 27 28 29 30 31 32 33 34 35 36 37 38 39
+ DPT_PCB3_1MHz_half
XY1 27 28 29 30 31 32 33 34 35 36 37 38 39 DPT_PCB3_1MHz_parlel
XZhalf2 27 28 29 30 31 32 33 34 35 36 37 38 39 14 14 14 15 16 16 17 18 19 20 20
+ 20 21 DPT_PCB3_1MHz_half

.subckt DPT_PCB3_1MHz_half 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21
+ 22 23 24 25 26
V1 1 27 dc 0.0
V2 2 28 dc 0.0
V3 3 29 dc 0.0
V4 4 30 dc 0.0
V5 5 31 dc 0.0
V6 6 32 dc 0.0
V7 7 33 dc 0.0
V8 8 34 dc 0.0
V9 9 35 dc 0.0
V10 10 36 dc 0.0
V11 11 37 dc 0.0
V12 12 38 dc 0.0
V13 13 39 dc 0.0
R1 27 40 0.0047064192961
R2 28 41 0.00695101712772
R3 29 42 0.00553905997109
R4 30 43 0.00387091111559
R5 31 44 0.00461604471545
R6 32 45 0.00693425524597
R7 33 46 0.00226380744624
R8 34 47 0.00452703279938
R9 35 48 0.00489886354568
R10 36 49 0.0138590154488
R11 37 50 0.0103844780021
R12 38 51 0.0185858928865
R13 39 52 0.00396873572192
F1_2 40 27 V2 0.510994
F1_3 40 27 V3 0.976857
F1_4 40 27 V4 -0.00664462
F1_5 40 27 V5 0.0213108
F1_6 40 27 V6 0.00956853
F1_7 40 27 V7 -0.0195748
F1_8 40 27 V8 0.0183497
F1_9 40 27 V9 -0.00598432
F1_10 40 27 V10 0.0881422
F1_11 40 27 V11 -0.0252051
F1_12 40 27 V12 -0.000938995
F1_13 40 27 V13 0.00308048
F2_1 41 28 V1 0.345985
F2_3 41 28 V3 0.345038
F2_4 41 28 V4 -0.00250735
F2_5 41 28 V5 0.00123936
F2_6 41 28 V6 -0.0102022
F2_7 41 28 V7 -0.00637351
F2_8 41 28 V8 0.0124154
F2_9 41 28 V9 -0.00189189
F2_10 41 28 V10 0.0154634
F2_11 41 28 V11 -0.00826472
F2_12 41 28 V12 0.00447951
F2_13 41 28 V13 1.63612e-05
F3_1 42 29 V1 0.830014
F3_2 42 29 V2 0.432991
F3_4 42 29 V4 -0.00659127
F3_5 42 29 V5 0.0239857
F3_6 42 29 V6 0.00698749
F3_7 42 29 V7 -0.00819215
F3_8 42 29 V8 0.0199576
F3_9 42 29 V9 -0.00569155
F3_10 42 29 V10 0.0335231
F3_11 42 29 V11 0.0496
F3_12 42 29 V12 0.0775213
F3_13 42 29 V13 0.000199033
F4_1 43 30 V1 -0.00807881
F4_2 43 30 V2 -0.00450246
F4_3 43 30 V3 -0.00943175
F4_5 43 30 V5 -0.00801277
F4_6 43 30 V6 -0.0086714
F4_7 43 30 V7 0.0226837
F4_8 43 30 V8 -0.00391422
F4_9 43 30 V9 0.0141197
F4_10 43 30 V10 -0.00496125
F4_11 43 30 V11 -0.0079672
F4_12 43 30 V12 -0.0163027
F4_13 43 30 V13 -0.0322311
F5_1 44 31 V1 0.021728
F5_2 44 31 V2 0.00186628
F5_3 44 31 V3 0.0287818
F5_4 44 31 V4 -0.00671933
F5_6 44 31 V6 1.0291
F5_7 44 31 V7 -0.0135043
F5_8 44 31 V8 0.0148228
F5_9 44 31 V9 -0.00540601
F5_10 44 31 V10 0.0285475
F5_11 44 31 V11 -0.0149683
F5_12 44 31 V12 -0.0011018
F5_13 44 31 V13 0.0021595
F6_1 45 32 V1 0.00649435
F6_2 45 32 V2 -0.0102269
F6_3 45 32 V3 0.00558158
F6_4 45 32 V4 -0.00484064
F6_5 45 32 V5 0.685057
F6_7 45 32 V7 -0.00638185
F6_8 45 32 V8 0.00879152
F6_9 45 32 V9 -0.00225505
F6_10 45 32 V10 0.0158636
F6_11 45 32 V11 -0.0182896
F6_12 45 32 V12 -0.0043827
F6_13 45 32 V13 5.44738e-05
F7_1 46 33 V1 -0.0406958
F7_2 46 33 V2 -0.0195698
F7_3 46 33 V3 -0.0200445
F7_4 46 33 V4 0.0387871
F7_5 46 33 V5 -0.0275361
F7_6 46 33 V6 -0.0195482
F7_8 46 33 V8 -0.0194336
F7_9 46 33 V9 0.0427568
F7_10 46 33 V10 -0.0364709
F7_11 46 33 V11 -0.128571
F7_12 46 33 V12 -0.23228
F7_13 46 33 V13 -0.0607442
F8_1 47 34 V1 0.0190768
F8_2 47 34 V2 0.0190631
F8_3 47 34 V3 0.0244192
F8_4 47 34 V4 -0.00334691
F8_5 47 34 V5 0.0151143
F8_6 47 34 V6 0.0134664
F8_7 47 34 V7 -0.00971805
F8_9 47 34 V9 -0.007398
F8_10 47 34 V10 0.0318493
F8_11 47 34 V11 0.0349783
F8_12 47 34 V12 0.0855572
F8_13 47 34 V13 0.00229397
F9_1 48 35 V1 -0.00574923
F9_2 48 35 V2 -0.00268441
F9_3 48 35 V3 -0.00643534
F9_4 48 35 V4 0.0111569
F9_5 48 35 V5 -0.00509392
F9_6 48 35 V6 -0.00319199
F9_7 48 35 V7 0.0197583
F9_8 48 35 V8 -0.00683648
F9_10 48 35 V10 -0.00414847
F9_11 48 35 V11 -0.0263781
F9_12 48 35 V12 -0.0338538
F9_13 48 35 V13 -0.00900641
F10_1 49 36 V1 0.0299325
F10_2 49 36 V2 0.0077557
F10_3 49 36 V3 0.0133983
F10_4 49 36 V4 -0.00138571
F10_5 49 36 V5 0.00950835
F10_6 49 36 V6 0.00793724
F10_7 49 36 V7 -0.00595735
F10_8 49 36 V8 0.0104035
F10_9 49 36 V9 -0.0014664
F10_11 49 36 V11 0.0303868
F10_12 49 36 V12 0.0410802
F10_13 49 36 V13 -0.000733903
F11_1 50 37 V1 -0.0114234
F11_2 50 37 V2 -0.00553213
F11_3 50 37 V3 0.0264566
F11_4 50 37 V4 -0.00296985
F11_5 50 37 V5 -0.00665363
F11_6 50 37 V6 -0.0122129
F11_7 50 37 V7 -0.0280284
F11_8 50 37 V8 0.0152485
F11_9 50 37 V9 -0.0124438
F11_10 50 37 V10 0.0405539
F11_12 50 37 V12 1.00422
F11_13 50 37 V13 0.00821434
F12_1 51 38 V1 -0.000237777
F12_2 51 38 V2 0.00167531
F12_3 51 38 V3 0.0231033
F12_4 51 38 V4 -0.00339539
F12_5 51 38 V5 -0.000273646
F12_6 51 38 V6 -0.00163515
F12_7 51 38 V7 -0.0282923
F12_8 51 38 V8 0.0208395
F12_9 51 38 V9 -0.00892317
F12_10 51 38 V10 0.0306324
F12_11 51 38 V11 0.561085
F12_13 51 38 V13 0.00581952
F13_1 52 39 V1 0.00365306
F13_2 52 39 V2 2.86556e-05
F13_3 52 39 V3 0.000277785
F13_4 52 39 V4 -0.0314366
F13_5 52 39 V5 0.00251172
F13_6 52 39 V6 9.51777e-05
F13_7 52 39 V7 -0.0346491
F13_8 52 39 V8 0.00261667
F13_9 52 39 V9 -0.0111172
F13_10 52 39 V10 -0.00256283
F13_11 52 39 V11 0.0214934
F13_12 52 39 V12 0.0272532
L1 40 14 1.36222321603e-08
L2 41 15 6.74519834081e-09
L3 42 16 1.48593610162e-08
L4 43 17 1.12776182766e-09
L5 44 18 8.20681777212e-09
L6 45 19 8.67829102419e-09
L7 46 20 1.751645696e-09
L8 47 21 3.33221255608e-09
L9 48 22 1.7551676085e-09
L10 49 23 1.10822348259e-08
L11 50 24 7.26259197051e-09
L12 51 25 1.21071860569e-08
L13 52 26 1.19932180095e-09
K1_2 L1 L2 0.570956
K1_3 L1 L3 0.926577
K1_4 L1 L4 -0.0148986
K1_5 L1 L5 0.0665765
K1_6 L1 L6 0.0547754
K1_7 L1 L7 -0.0296063
K1_8 L1 L8 0.0207254
K1_9 L1 L9 -0.00998227
K1_10 L1 L10 0.073468
K1_11 L1 L11 -0.00750816
K1_12 L1 L12 0.0156907
K1_13 L1 L13 0.00437073
K2_3 L2 L3 0.544393
K2_4 L2 L4 -0.00824377
K2_5 L2 L5 0.0565616
K2_6 L2 L6 0.0465712
K2_7 L2 L7 -0.0151074
K2_8 L2 L8 0.0117472
K2_9 L2 L9 -0.00480209
K2_10 L2 L10 0.0247228
K2_11 L2 L11 -0.00537154
K2_12 L2 L12 0.00671203
K2_13 L2 L13 0.00161785
K3_4 L3 L4 -0.0157076
K3_5 L3 L5 0.0677713
K3_6 L3 L6 0.0559359
K3_7 L3 L7 -0.0316337
K3_8 L3 L8 0.0220344
K3_9 L3 L9 -0.0137088
K3_10 L3 L10 0.0132005
K3_11 L3 L11 0.0244726
K3_12 L3 L12 0.0400461
K3_13 L3 L13 0.00707002
K4_5 L4 L5 -0.0172219
K4_6 L4 L6 -0.0154487
K4_7 L4 L7 0.0899754
K4_8 L4 L8 -0.0130395
K4_9 L4 L9 0.0243238
K4_10 L4 L10 -0.00878857
K4_11 L4 L11 -0.00041469
K4_12 L4 L12 -0.0285952
K4_13 L4 L13 -0.179574
K5_6 L5 L6 0.945712
K5_7 L5 L7 -0.0334898
K5_8 L5 L8 0.018975
K5_9 L5 L9 -0.0141429
K5_10 L5 L10 0.0131524
K5_11 L5 L11 0.00129649
K5_12 L5 L12 0.0170612
K5_13 L5 L13 0.00824276
K6_7 L6 L7 -0.0292692
K6_8 L6 L8 0.014891
K6_9 L6 L9 -0.0123744
K6_10 L6 L10 0.0106018
K6_11 L6 L11 0.00066583
K6_12 L6 L12 0.0147578
K6_13 L6 L13 0.00732007
K7_8 L7 L8 -0.0422198
K7_9 L7 L9 0.330245
K7_10 L7 L10 -0.012784
K7_11 L7 L11 -0.0261832
K7_12 L7 L12 -0.145188
K7_13 L7 L13 -0.0723898
K8_9 L8 L9 -0.0268091
K8_10 L8 L10 0.0105446
K8_11 L8 L11 0.0128639
K8_12 L8 L12 0.0399591
K8_13 L8 L13 0.00699401
K9_10 L9 L10 -0.00170648
K9_11 L9 L11 -0.017482
K9_12 L9 L12 -0.0619707
K9_13 L9 L13 -0.0371575
K10_11 L10 L11 -0.00964367
K10_12 L10 L12 0.0113708
K10_13 L10 L13 -0.00150318
K11_12 L11 L12 0.76148
K11_13 L11 L13 0.01251
K12_13 L12 L13 0.0245034
.ends DPT_PCB3_1MHz_half

.subckt DPT_PCB3_1MHz_parlel 1 2 3 4 5 6 7 8 9 10 11 12 13
RG1_4 1 4 784315927990
RG1_5 1 5 101236329.706
RG1_6 1 6 101236329.706
RG1_7 1 7 -5234806651.55
RG1_8 1 8 1616629975.37
RG1_9 1 9 -463085456175
RG1_10 1 10 943903488.117
RG1_11 1 11 943903488.117
RG1_12 1 12 943903488.117
RG1_13 1 13 -554400132949
RG2_4 2 4 784315927990
RG2_5 2 5 101236329.706
RG2_6 2 6 101236329.706
RG2_7 2 7 -5234806651.55
RG2_8 2 8 1616629975.37
RG2_9 2 9 -463085456175
RG2_10 2 10 943903488.117
RG2_11 2 11 943903488.117
RG2_12 2 12 943903488.117
RG2_13 2 13 -554400132949
RG3_4 3 4 784315927990
RG3_5 3 5 101236329.706
RG3_6 3 6 101236329.706
RG3_7 3 7 -5234806651.55
RG3_8 3 8 1616629975.37
RG3_9 3 9 -463085456175
RG3_10 3 10 943903488.117
RG3_11 3 11 943903488.117
RG3_12 3 12 943903488.117
RG3_13 3 13 -554400132949
R4_0 4 0 22778316.9718
RG4_5 4 5 -92955802664
RG4_6 4 6 -92955802664
RG4_7 4 7 229932185.722
RG4_8 4 8 991387515865
RG4_9 4 9 -131136135670
RG4_10 4 10 -936757114203
RG4_11 4 11 -936757114203
RG4_12 4 12 -936757114203
RG4_13 4 13 63044174.374
RG5_7 5 7 2220831416.18
RG5_8 5 8 63238135.3782
RG5_9 5 9 -21290853316.3
RG5_10 5 10 35247616685.5
RG5_11 5 11 35247616685.5
RG5_12 5 12 35247616685.5
RG5_13 5 13 -27357990048.5
RG6_7 6 7 2220831416.18
RG6_8 6 8 63238135.3782
RG6_9 6 9 -21290853316.3
RG6_10 6 10 35247616685.5
RG6_11 6 11 35247616685.5
RG6_12 6 12 35247616685.5
RG6_13 6 13 -27357990048.5
R7_0 7 0 2618210.82461
RG7_8 7 8 42796515.7764
RG7_9 7 9 4198671.78536
RG7_10 7 10 99576611.9066
RG7_11 7 11 99576611.9066
RG7_12 7 12 99576611.9066
RG7_13 7 13 6776230.8102
R8_0 8 0 433126698.518
RG8_9 8 9 -15297776473.2
RG8_10 8 10 687288198.303
RG8_11 8 11 687288198.303
RG8_12 8 12 687288198.303
RG8_13 8 13 -191138532056
RG9_10 9 10 1.10220470938e+12
RG9_11 9 11 1.10220470938e+12
RG9_12 9 12 1.10220470938e+12
RG9_13 9 13 -383976657399
R10_0 10 0 165180165.963
RG10_13 10 13 -178965163267
R11_0 11 0 165180165.963
RG11_13 11 13 -178965163267
R12_0 12 0 165180165.963
RG12_13 12 13 -178965163267
R13_0 13 0 175782103.272
C1_0 1 0 5.0578024213e-13
C1_4 1 4 7.67944644702e-17
C1_5 1 5 4.56160147835e-13
C1_6 1 6 4.56160147835e-13
C1_7 1 7 1.23782970253e-13
C1_8 1 8 6.40385295255e-14
C1_9 1 9 6.76056100866e-16
C1_10 1 10 4.05813908766e-14
C1_11 1 11 4.05813908766e-14
C1_12 1 12 4.05813908766e-14
C1_13 1 13 1.13444400204e-15
C2_0 2 0 5.0578024213e-13
C2_4 2 4 7.67944644702e-17
C2_5 2 5 4.56160147835e-13
C2_6 2 6 4.56160147835e-13
C2_7 2 7 1.23782970253e-13
C2_8 2 8 6.40385295255e-14
C2_9 2 9 6.76056100866e-16
C2_10 2 10 4.05813908766e-14
C2_11 2 11 4.05813908766e-14
C2_12 2 12 4.05813908766e-14
C2_13 2 13 1.13444400204e-15
C3_0 3 0 5.0578024213e-13
C3_4 3 4 7.67944644702e-17
C3_5 3 5 4.56160147835e-13
C3_6 3 6 4.56160147835e-13
C3_7 3 7 1.23782970253e-13
C3_8 3 8 6.40385295255e-14
C3_9 3 9 6.76056100866e-16
C3_10 3 10 4.05813908766e-14
C3_11 3 11 4.05813908766e-14
C3_12 3 12 4.05813908766e-14
C3_13 3 13 1.13444400204e-15
C4_0 4 0 4.46914732367e-13
C4_5 4 5 1.15696949489e-16
C4_6 4 6 1.15696949489e-16
C4_7 4 7 7.30852207514e-14
C4_8 4 8 2.44789613597e-16
C4_9 4 9 1.37905258181e-16
C4_10 4 10 4.68211949804e-17
C4_11 4 11 4.68211949804e-17
C4_12 4 12 4.68211949804e-17
C4_13 4 13 1.74165702734e-13
C5_0 5 0 7.10021301952e-13
C5_7 5 7 2.71661205128e-13
C5_8 5 8 5.28803675544e-13
C5_9 5 9 1.88203286195e-15
C5_10 5 10 8.92687168925e-15
C5_11 5 11 8.92687168925e-15
C5_12 5 12 8.92687168925e-15
C5_13 5 13 2.05581185292e-15
C6_0 6 0 7.10021301952e-13
C6_7 6 7 2.71661205128e-13
C6_8 6 8 5.28803675544e-13
C6_9 6 9 1.88203286195e-15
C6_10 6 10 8.92687168925e-15
C6_11 6 11 8.92687168925e-15
C6_12 6 12 8.92687168925e-15
C6_13 6 13 2.05581185292e-15
C7_0 7 0 5.89738570442e-12
C7_8 7 8 7.14624610461e-13
C7_9 7 9 2.58821852452e-12
C7_10 7 10 3.00272699964e-13
C7_11 7 11 3.00272699964e-13
C7_12 7 12 3.00272699964e-13
C7_13 7 13 2.33918218628e-12
C8_0 8 0 1.35172475367e-13
C8_9 8 9 1.03667900422e-14
C8_10 8 10 4.99628648661e-14
C8_11 8 11 4.99628648661e-14
C8_12 8 12 4.99628648661e-14
C8_13 8 13 1.93537057557e-15
C9_10 9 10 1.46824125633e-15
C9_11 9 11 1.46824125633e-15
C9_12 9 12 1.46824125633e-15
C9_13 9 13 7.27265029604e-16
C10_0 10 0 1.56201216817e-13
C10_13 10 13 9.12598687274e-16
C11_0 11 0 1.56201216817e-13
C11_13 11 13 9.12598687274e-16
C12_0 12 0 1.56201216817e-13
C12_13 12 13 9.12598687274e-16
C13_0 13 0 1.3169689766e-13
.ends DPT_PCB3_1MHz_parlel

.ends DPT_PCB3_1MHz
